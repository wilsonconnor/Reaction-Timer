module binaryToBCDRam(
    input clk,
    input [15:0] val,
    output reg [3:0] bcd3,
    output reg [3:0] bcd2,
    output reg [3:0] bcd1,
    output reg [3:0] bcd0
    );
    
    always@(posedge clk)
    begin
    case(val)
    
			0: begin bcd3<=0;bcd2<=0;bcd1<=0;bcd0<=0; end
			1: begin bcd3<=0;bcd2<=0;bcd1<=0;bcd0<=1; end
			2: begin bcd3<=0;bcd2<=0;bcd1<=0;bcd0<=2; end
			3: begin bcd3<=0;bcd2<=0;bcd1<=0;bcd0<=3; end
			4: begin bcd3<=0;bcd2<=0;bcd1<=0;bcd0<=4; end
			5: begin bcd3<=0;bcd2<=0;bcd1<=0;bcd0<=5; end
			6: begin bcd3<=0;bcd2<=0;bcd1<=0;bcd0<=6; end
			7: begin bcd3<=0;bcd2<=0;bcd1<=0;bcd0<=7; end
			8: begin bcd3<=0;bcd2<=0;bcd1<=0;bcd0<=8; end
			9: begin bcd3<=0;bcd2<=0;bcd1<=0;bcd0<=9; end
			10: begin bcd3<=0;bcd2<=0;bcd1<=1;bcd0<=0; end
			11: begin bcd3<=0;bcd2<=0;bcd1<=1;bcd0<=1; end
			12: begin bcd3<=0;bcd2<=0;bcd1<=1;bcd0<=2; end
			13: begin bcd3<=0;bcd2<=0;bcd1<=1;bcd0<=3; end
			14: begin bcd3<=0;bcd2<=0;bcd1<=1;bcd0<=4; end
			15: begin bcd3<=0;bcd2<=0;bcd1<=1;bcd0<=5; end
			16: begin bcd3<=0;bcd2<=0;bcd1<=1;bcd0<=6; end
			17: begin bcd3<=0;bcd2<=0;bcd1<=1;bcd0<=7; end
			18: begin bcd3<=0;bcd2<=0;bcd1<=1;bcd0<=8; end
			19: begin bcd3<=0;bcd2<=0;bcd1<=1;bcd0<=9; end
			20: begin bcd3<=0;bcd2<=0;bcd1<=2;bcd0<=0; end
			21: begin bcd3<=0;bcd2<=0;bcd1<=2;bcd0<=1; end
			22: begin bcd3<=0;bcd2<=0;bcd1<=2;bcd0<=2; end
			23: begin bcd3<=0;bcd2<=0;bcd1<=2;bcd0<=3; end
			24: begin bcd3<=0;bcd2<=0;bcd1<=2;bcd0<=4; end
			25: begin bcd3<=0;bcd2<=0;bcd1<=2;bcd0<=5; end
			26: begin bcd3<=0;bcd2<=0;bcd1<=2;bcd0<=6; end
			27: begin bcd3<=0;bcd2<=0;bcd1<=2;bcd0<=7; end
			28: begin bcd3<=0;bcd2<=0;bcd1<=2;bcd0<=8; end
			29: begin bcd3<=0;bcd2<=0;bcd1<=2;bcd0<=9; end
			30: begin bcd3<=0;bcd2<=0;bcd1<=3;bcd0<=0; end
			31: begin bcd3<=0;bcd2<=0;bcd1<=3;bcd0<=1; end
			32: begin bcd3<=0;bcd2<=0;bcd1<=3;bcd0<=2; end
			33: begin bcd3<=0;bcd2<=0;bcd1<=3;bcd0<=3; end
			34: begin bcd3<=0;bcd2<=0;bcd1<=3;bcd0<=4; end
			35: begin bcd3<=0;bcd2<=0;bcd1<=3;bcd0<=5; end
			36: begin bcd3<=0;bcd2<=0;bcd1<=3;bcd0<=6; end
			37: begin bcd3<=0;bcd2<=0;bcd1<=3;bcd0<=7; end
			38: begin bcd3<=0;bcd2<=0;bcd1<=3;bcd0<=8; end
			39: begin bcd3<=0;bcd2<=0;bcd1<=3;bcd0<=9; end
			40: begin bcd3<=0;bcd2<=0;bcd1<=4;bcd0<=0; end
			41: begin bcd3<=0;bcd2<=0;bcd1<=4;bcd0<=1; end
			42: begin bcd3<=0;bcd2<=0;bcd1<=4;bcd0<=2; end
			43: begin bcd3<=0;bcd2<=0;bcd1<=4;bcd0<=3; end
			44: begin bcd3<=0;bcd2<=0;bcd1<=4;bcd0<=4; end
			45: begin bcd3<=0;bcd2<=0;bcd1<=4;bcd0<=5; end
			46: begin bcd3<=0;bcd2<=0;bcd1<=4;bcd0<=6; end
			47: begin bcd3<=0;bcd2<=0;bcd1<=4;bcd0<=7; end
			48: begin bcd3<=0;bcd2<=0;bcd1<=4;bcd0<=8; end
			49: begin bcd3<=0;bcd2<=0;bcd1<=4;bcd0<=9; end
			50: begin bcd3<=0;bcd2<=0;bcd1<=5;bcd0<=0; end
			51: begin bcd3<=0;bcd2<=0;bcd1<=5;bcd0<=1; end
			52: begin bcd3<=0;bcd2<=0;bcd1<=5;bcd0<=2; end
			53: begin bcd3<=0;bcd2<=0;bcd1<=5;bcd0<=3; end
			54: begin bcd3<=0;bcd2<=0;bcd1<=5;bcd0<=4; end
			55: begin bcd3<=0;bcd2<=0;bcd1<=5;bcd0<=5; end
			56: begin bcd3<=0;bcd2<=0;bcd1<=5;bcd0<=6; end
			57: begin bcd3<=0;bcd2<=0;bcd1<=5;bcd0<=7; end
			58: begin bcd3<=0;bcd2<=0;bcd1<=5;bcd0<=8; end
			59: begin bcd3<=0;bcd2<=0;bcd1<=5;bcd0<=9; end
			60: begin bcd3<=0;bcd2<=0;bcd1<=6;bcd0<=0; end
			61: begin bcd3<=0;bcd2<=0;bcd1<=6;bcd0<=1; end
			62: begin bcd3<=0;bcd2<=0;bcd1<=6;bcd0<=2; end
			63: begin bcd3<=0;bcd2<=0;bcd1<=6;bcd0<=3; end
			64: begin bcd3<=0;bcd2<=0;bcd1<=6;bcd0<=4; end
			65: begin bcd3<=0;bcd2<=0;bcd1<=6;bcd0<=5; end
			66: begin bcd3<=0;bcd2<=0;bcd1<=6;bcd0<=6; end
			67: begin bcd3<=0;bcd2<=0;bcd1<=6;bcd0<=7; end
			68: begin bcd3<=0;bcd2<=0;bcd1<=6;bcd0<=8; end
			69: begin bcd3<=0;bcd2<=0;bcd1<=6;bcd0<=9; end
			70: begin bcd3<=0;bcd2<=0;bcd1<=7;bcd0<=0; end
			71: begin bcd3<=0;bcd2<=0;bcd1<=7;bcd0<=1; end
			72: begin bcd3<=0;bcd2<=0;bcd1<=7;bcd0<=2; end
			73: begin bcd3<=0;bcd2<=0;bcd1<=7;bcd0<=3; end
			74: begin bcd3<=0;bcd2<=0;bcd1<=7;bcd0<=4; end
			75: begin bcd3<=0;bcd2<=0;bcd1<=7;bcd0<=5; end
			76: begin bcd3<=0;bcd2<=0;bcd1<=7;bcd0<=6; end
			77: begin bcd3<=0;bcd2<=0;bcd1<=7;bcd0<=7; end
			78: begin bcd3<=0;bcd2<=0;bcd1<=7;bcd0<=8; end
			79: begin bcd3<=0;bcd2<=0;bcd1<=7;bcd0<=9; end
			80: begin bcd3<=0;bcd2<=0;bcd1<=8;bcd0<=0; end
			81: begin bcd3<=0;bcd2<=0;bcd1<=8;bcd0<=1; end
			82: begin bcd3<=0;bcd2<=0;bcd1<=8;bcd0<=2; end
			83: begin bcd3<=0;bcd2<=0;bcd1<=8;bcd0<=3; end
			84: begin bcd3<=0;bcd2<=0;bcd1<=8;bcd0<=4; end
			85: begin bcd3<=0;bcd2<=0;bcd1<=8;bcd0<=5; end
			86: begin bcd3<=0;bcd2<=0;bcd1<=8;bcd0<=6; end
			87: begin bcd3<=0;bcd2<=0;bcd1<=8;bcd0<=7; end
			88: begin bcd3<=0;bcd2<=0;bcd1<=8;bcd0<=8; end
			89: begin bcd3<=0;bcd2<=0;bcd1<=8;bcd0<=9; end
			90: begin bcd3<=0;bcd2<=0;bcd1<=9;bcd0<=0; end
			91: begin bcd3<=0;bcd2<=0;bcd1<=9;bcd0<=1; end
			92: begin bcd3<=0;bcd2<=0;bcd1<=9;bcd0<=2; end
			93: begin bcd3<=0;bcd2<=0;bcd1<=9;bcd0<=3; end
			94: begin bcd3<=0;bcd2<=0;bcd1<=9;bcd0<=4; end
			95: begin bcd3<=0;bcd2<=0;bcd1<=9;bcd0<=5; end
			96: begin bcd3<=0;bcd2<=0;bcd1<=9;bcd0<=6; end
			97: begin bcd3<=0;bcd2<=0;bcd1<=9;bcd0<=7; end
			98: begin bcd3<=0;bcd2<=0;bcd1<=9;bcd0<=8; end
			99: begin bcd3<=0;bcd2<=0;bcd1<=9;bcd0<=9; end
			100: begin bcd3<=0;bcd2<=1;bcd1<=0;bcd0<=0; end
			101: begin bcd3<=0;bcd2<=1;bcd1<=0;bcd0<=1; end
			102: begin bcd3<=0;bcd2<=1;bcd1<=0;bcd0<=2; end
			103: begin bcd3<=0;bcd2<=1;bcd1<=0;bcd0<=3; end
			104: begin bcd3<=0;bcd2<=1;bcd1<=0;bcd0<=4; end
			105: begin bcd3<=0;bcd2<=1;bcd1<=0;bcd0<=5; end
			106: begin bcd3<=0;bcd2<=1;bcd1<=0;bcd0<=6; end
			107: begin bcd3<=0;bcd2<=1;bcd1<=0;bcd0<=7; end
			108: begin bcd3<=0;bcd2<=1;bcd1<=0;bcd0<=8; end
			109: begin bcd3<=0;bcd2<=1;bcd1<=0;bcd0<=9; end
			110: begin bcd3<=0;bcd2<=1;bcd1<=1;bcd0<=0; end
			111: begin bcd3<=0;bcd2<=1;bcd1<=1;bcd0<=1; end
			112: begin bcd3<=0;bcd2<=1;bcd1<=1;bcd0<=2; end
			113: begin bcd3<=0;bcd2<=1;bcd1<=1;bcd0<=3; end
			114: begin bcd3<=0;bcd2<=1;bcd1<=1;bcd0<=4; end
			115: begin bcd3<=0;bcd2<=1;bcd1<=1;bcd0<=5; end
			116: begin bcd3<=0;bcd2<=1;bcd1<=1;bcd0<=6; end
			117: begin bcd3<=0;bcd2<=1;bcd1<=1;bcd0<=7; end
			118: begin bcd3<=0;bcd2<=1;bcd1<=1;bcd0<=8; end
			119: begin bcd3<=0;bcd2<=1;bcd1<=1;bcd0<=9; end
			120: begin bcd3<=0;bcd2<=1;bcd1<=2;bcd0<=0; end
			121: begin bcd3<=0;bcd2<=1;bcd1<=2;bcd0<=1; end
			122: begin bcd3<=0;bcd2<=1;bcd1<=2;bcd0<=2; end
			123: begin bcd3<=0;bcd2<=1;bcd1<=2;bcd0<=3; end
			124: begin bcd3<=0;bcd2<=1;bcd1<=2;bcd0<=4; end
			125: begin bcd3<=0;bcd2<=1;bcd1<=2;bcd0<=5; end
			126: begin bcd3<=0;bcd2<=1;bcd1<=2;bcd0<=6; end
			127: begin bcd3<=0;bcd2<=1;bcd1<=2;bcd0<=7; end
			128: begin bcd3<=0;bcd2<=1;bcd1<=2;bcd0<=8; end
			129: begin bcd3<=0;bcd2<=1;bcd1<=2;bcd0<=9; end
			130: begin bcd3<=0;bcd2<=1;bcd1<=3;bcd0<=0; end
			131: begin bcd3<=0;bcd2<=1;bcd1<=3;bcd0<=1; end
			132: begin bcd3<=0;bcd2<=1;bcd1<=3;bcd0<=2; end
			133: begin bcd3<=0;bcd2<=1;bcd1<=3;bcd0<=3; end
			134: begin bcd3<=0;bcd2<=1;bcd1<=3;bcd0<=4; end
			135: begin bcd3<=0;bcd2<=1;bcd1<=3;bcd0<=5; end
			136: begin bcd3<=0;bcd2<=1;bcd1<=3;bcd0<=6; end
			137: begin bcd3<=0;bcd2<=1;bcd1<=3;bcd0<=7; end
			138: begin bcd3<=0;bcd2<=1;bcd1<=3;bcd0<=8; end
			139: begin bcd3<=0;bcd2<=1;bcd1<=3;bcd0<=9; end
			140: begin bcd3<=0;bcd2<=1;bcd1<=4;bcd0<=0; end
			141: begin bcd3<=0;bcd2<=1;bcd1<=4;bcd0<=1; end
			142: begin bcd3<=0;bcd2<=1;bcd1<=4;bcd0<=2; end
			143: begin bcd3<=0;bcd2<=1;bcd1<=4;bcd0<=3; end
			144: begin bcd3<=0;bcd2<=1;bcd1<=4;bcd0<=4; end
			145: begin bcd3<=0;bcd2<=1;bcd1<=4;bcd0<=5; end
			146: begin bcd3<=0;bcd2<=1;bcd1<=4;bcd0<=6; end
			147: begin bcd3<=0;bcd2<=1;bcd1<=4;bcd0<=7; end
			148: begin bcd3<=0;bcd2<=1;bcd1<=4;bcd0<=8; end
			149: begin bcd3<=0;bcd2<=1;bcd1<=4;bcd0<=9; end
			150: begin bcd3<=0;bcd2<=1;bcd1<=5;bcd0<=0; end
			151: begin bcd3<=0;bcd2<=1;bcd1<=5;bcd0<=1; end
			152: begin bcd3<=0;bcd2<=1;bcd1<=5;bcd0<=2; end
			153: begin bcd3<=0;bcd2<=1;bcd1<=5;bcd0<=3; end
			154: begin bcd3<=0;bcd2<=1;bcd1<=5;bcd0<=4; end
			155: begin bcd3<=0;bcd2<=1;bcd1<=5;bcd0<=5; end
			156: begin bcd3<=0;bcd2<=1;bcd1<=5;bcd0<=6; end
			157: begin bcd3<=0;bcd2<=1;bcd1<=5;bcd0<=7; end
			158: begin bcd3<=0;bcd2<=1;bcd1<=5;bcd0<=8; end
			159: begin bcd3<=0;bcd2<=1;bcd1<=5;bcd0<=9; end
			160: begin bcd3<=0;bcd2<=1;bcd1<=6;bcd0<=0; end
			161: begin bcd3<=0;bcd2<=1;bcd1<=6;bcd0<=1; end
			162: begin bcd3<=0;bcd2<=1;bcd1<=6;bcd0<=2; end
			163: begin bcd3<=0;bcd2<=1;bcd1<=6;bcd0<=3; end
			164: begin bcd3<=0;bcd2<=1;bcd1<=6;bcd0<=4; end
			165: begin bcd3<=0;bcd2<=1;bcd1<=6;bcd0<=5; end
			166: begin bcd3<=0;bcd2<=1;bcd1<=6;bcd0<=6; end
			167: begin bcd3<=0;bcd2<=1;bcd1<=6;bcd0<=7; end
			168: begin bcd3<=0;bcd2<=1;bcd1<=6;bcd0<=8; end
			169: begin bcd3<=0;bcd2<=1;bcd1<=6;bcd0<=9; end
			170: begin bcd3<=0;bcd2<=1;bcd1<=7;bcd0<=0; end
			171: begin bcd3<=0;bcd2<=1;bcd1<=7;bcd0<=1; end
			172: begin bcd3<=0;bcd2<=1;bcd1<=7;bcd0<=2; end
			173: begin bcd3<=0;bcd2<=1;bcd1<=7;bcd0<=3; end
			174: begin bcd3<=0;bcd2<=1;bcd1<=7;bcd0<=4; end
			175: begin bcd3<=0;bcd2<=1;bcd1<=7;bcd0<=5; end
			176: begin bcd3<=0;bcd2<=1;bcd1<=7;bcd0<=6; end
			177: begin bcd3<=0;bcd2<=1;bcd1<=7;bcd0<=7; end
			178: begin bcd3<=0;bcd2<=1;bcd1<=7;bcd0<=8; end
			179: begin bcd3<=0;bcd2<=1;bcd1<=7;bcd0<=9; end
			180: begin bcd3<=0;bcd2<=1;bcd1<=8;bcd0<=0; end
			181: begin bcd3<=0;bcd2<=1;bcd1<=8;bcd0<=1; end
			182: begin bcd3<=0;bcd2<=1;bcd1<=8;bcd0<=2; end
			183: begin bcd3<=0;bcd2<=1;bcd1<=8;bcd0<=3; end
			184: begin bcd3<=0;bcd2<=1;bcd1<=8;bcd0<=4; end
			185: begin bcd3<=0;bcd2<=1;bcd1<=8;bcd0<=5; end
			186: begin bcd3<=0;bcd2<=1;bcd1<=8;bcd0<=6; end
			187: begin bcd3<=0;bcd2<=1;bcd1<=8;bcd0<=7; end
			188: begin bcd3<=0;bcd2<=1;bcd1<=8;bcd0<=8; end
			189: begin bcd3<=0;bcd2<=1;bcd1<=8;bcd0<=9; end
			190: begin bcd3<=0;bcd2<=1;bcd1<=9;bcd0<=0; end
			191: begin bcd3<=0;bcd2<=1;bcd1<=9;bcd0<=1; end
			192: begin bcd3<=0;bcd2<=1;bcd1<=9;bcd0<=2; end
			193: begin bcd3<=0;bcd2<=1;bcd1<=9;bcd0<=3; end
			194: begin bcd3<=0;bcd2<=1;bcd1<=9;bcd0<=4; end
			195: begin bcd3<=0;bcd2<=1;bcd1<=9;bcd0<=5; end
			196: begin bcd3<=0;bcd2<=1;bcd1<=9;bcd0<=6; end
			197: begin bcd3<=0;bcd2<=1;bcd1<=9;bcd0<=7; end
			198: begin bcd3<=0;bcd2<=1;bcd1<=9;bcd0<=8; end
			199: begin bcd3<=0;bcd2<=1;bcd1<=9;bcd0<=9; end
			200: begin bcd3<=0;bcd2<=2;bcd1<=0;bcd0<=0; end
			201: begin bcd3<=0;bcd2<=2;bcd1<=0;bcd0<=1; end
			202: begin bcd3<=0;bcd2<=2;bcd1<=0;bcd0<=2; end
			203: begin bcd3<=0;bcd2<=2;bcd1<=0;bcd0<=3; end
			204: begin bcd3<=0;bcd2<=2;bcd1<=0;bcd0<=4; end
			205: begin bcd3<=0;bcd2<=2;bcd1<=0;bcd0<=5; end
			206: begin bcd3<=0;bcd2<=2;bcd1<=0;bcd0<=6; end
			207: begin bcd3<=0;bcd2<=2;bcd1<=0;bcd0<=7; end
			208: begin bcd3<=0;bcd2<=2;bcd1<=0;bcd0<=8; end
			209: begin bcd3<=0;bcd2<=2;bcd1<=0;bcd0<=9; end
			210: begin bcd3<=0;bcd2<=2;bcd1<=1;bcd0<=0; end
			211: begin bcd3<=0;bcd2<=2;bcd1<=1;bcd0<=1; end
			212: begin bcd3<=0;bcd2<=2;bcd1<=1;bcd0<=2; end
			213: begin bcd3<=0;bcd2<=2;bcd1<=1;bcd0<=3; end
			214: begin bcd3<=0;bcd2<=2;bcd1<=1;bcd0<=4; end
			215: begin bcd3<=0;bcd2<=2;bcd1<=1;bcd0<=5; end
			216: begin bcd3<=0;bcd2<=2;bcd1<=1;bcd0<=6; end
			217: begin bcd3<=0;bcd2<=2;bcd1<=1;bcd0<=7; end
			218: begin bcd3<=0;bcd2<=2;bcd1<=1;bcd0<=8; end
			219: begin bcd3<=0;bcd2<=2;bcd1<=1;bcd0<=9; end
			220: begin bcd3<=0;bcd2<=2;bcd1<=2;bcd0<=0; end
			221: begin bcd3<=0;bcd2<=2;bcd1<=2;bcd0<=1; end
			222: begin bcd3<=0;bcd2<=2;bcd1<=2;bcd0<=2; end
			223: begin bcd3<=0;bcd2<=2;bcd1<=2;bcd0<=3; end
			224: begin bcd3<=0;bcd2<=2;bcd1<=2;bcd0<=4; end
			225: begin bcd3<=0;bcd2<=2;bcd1<=2;bcd0<=5; end
			226: begin bcd3<=0;bcd2<=2;bcd1<=2;bcd0<=6; end
			227: begin bcd3<=0;bcd2<=2;bcd1<=2;bcd0<=7; end
			228: begin bcd3<=0;bcd2<=2;bcd1<=2;bcd0<=8; end
			229: begin bcd3<=0;bcd2<=2;bcd1<=2;bcd0<=9; end
			230: begin bcd3<=0;bcd2<=2;bcd1<=3;bcd0<=0; end
			231: begin bcd3<=0;bcd2<=2;bcd1<=3;bcd0<=1; end
			232: begin bcd3<=0;bcd2<=2;bcd1<=3;bcd0<=2; end
			233: begin bcd3<=0;bcd2<=2;bcd1<=3;bcd0<=3; end
			234: begin bcd3<=0;bcd2<=2;bcd1<=3;bcd0<=4; end
			235: begin bcd3<=0;bcd2<=2;bcd1<=3;bcd0<=5; end
			236: begin bcd3<=0;bcd2<=2;bcd1<=3;bcd0<=6; end
			237: begin bcd3<=0;bcd2<=2;bcd1<=3;bcd0<=7; end
			238: begin bcd3<=0;bcd2<=2;bcd1<=3;bcd0<=8; end
			239: begin bcd3<=0;bcd2<=2;bcd1<=3;bcd0<=9; end
			240: begin bcd3<=0;bcd2<=2;bcd1<=4;bcd0<=0; end
			241: begin bcd3<=0;bcd2<=2;bcd1<=4;bcd0<=1; end
			242: begin bcd3<=0;bcd2<=2;bcd1<=4;bcd0<=2; end
			243: begin bcd3<=0;bcd2<=2;bcd1<=4;bcd0<=3; end
			244: begin bcd3<=0;bcd2<=2;bcd1<=4;bcd0<=4; end
			245: begin bcd3<=0;bcd2<=2;bcd1<=4;bcd0<=5; end
			246: begin bcd3<=0;bcd2<=2;bcd1<=4;bcd0<=6; end
			247: begin bcd3<=0;bcd2<=2;bcd1<=4;bcd0<=7; end
			248: begin bcd3<=0;bcd2<=2;bcd1<=4;bcd0<=8; end
			249: begin bcd3<=0;bcd2<=2;bcd1<=4;bcd0<=9; end
			250: begin bcd3<=0;bcd2<=2;bcd1<=5;bcd0<=0; end
			251: begin bcd3<=0;bcd2<=2;bcd1<=5;bcd0<=1; end
			252: begin bcd3<=0;bcd2<=2;bcd1<=5;bcd0<=2; end
			253: begin bcd3<=0;bcd2<=2;bcd1<=5;bcd0<=3; end
			254: begin bcd3<=0;bcd2<=2;bcd1<=5;bcd0<=4; end
			255: begin bcd3<=0;bcd2<=2;bcd1<=5;bcd0<=5; end
			256: begin bcd3<=0;bcd2<=2;bcd1<=5;bcd0<=6; end
			257: begin bcd3<=0;bcd2<=2;bcd1<=5;bcd0<=7; end
			258: begin bcd3<=0;bcd2<=2;bcd1<=5;bcd0<=8; end
			259: begin bcd3<=0;bcd2<=2;bcd1<=5;bcd0<=9; end
			260: begin bcd3<=0;bcd2<=2;bcd1<=6;bcd0<=0; end
			261: begin bcd3<=0;bcd2<=2;bcd1<=6;bcd0<=1; end
			262: begin bcd3<=0;bcd2<=2;bcd1<=6;bcd0<=2; end
			263: begin bcd3<=0;bcd2<=2;bcd1<=6;bcd0<=3; end
			264: begin bcd3<=0;bcd2<=2;bcd1<=6;bcd0<=4; end
			265: begin bcd3<=0;bcd2<=2;bcd1<=6;bcd0<=5; end
			266: begin bcd3<=0;bcd2<=2;bcd1<=6;bcd0<=6; end
			267: begin bcd3<=0;bcd2<=2;bcd1<=6;bcd0<=7; end
			268: begin bcd3<=0;bcd2<=2;bcd1<=6;bcd0<=8; end
			269: begin bcd3<=0;bcd2<=2;bcd1<=6;bcd0<=9; end
			270: begin bcd3<=0;bcd2<=2;bcd1<=7;bcd0<=0; end
			271: begin bcd3<=0;bcd2<=2;bcd1<=7;bcd0<=1; end
			272: begin bcd3<=0;bcd2<=2;bcd1<=7;bcd0<=2; end
			273: begin bcd3<=0;bcd2<=2;bcd1<=7;bcd0<=3; end
			274: begin bcd3<=0;bcd2<=2;bcd1<=7;bcd0<=4; end
			275: begin bcd3<=0;bcd2<=2;bcd1<=7;bcd0<=5; end
			276: begin bcd3<=0;bcd2<=2;bcd1<=7;bcd0<=6; end
			277: begin bcd3<=0;bcd2<=2;bcd1<=7;bcd0<=7; end
			278: begin bcd3<=0;bcd2<=2;bcd1<=7;bcd0<=8; end
			279: begin bcd3<=0;bcd2<=2;bcd1<=7;bcd0<=9; end
			280: begin bcd3<=0;bcd2<=2;bcd1<=8;bcd0<=0; end
			281: begin bcd3<=0;bcd2<=2;bcd1<=8;bcd0<=1; end
			282: begin bcd3<=0;bcd2<=2;bcd1<=8;bcd0<=2; end
			283: begin bcd3<=0;bcd2<=2;bcd1<=8;bcd0<=3; end
			284: begin bcd3<=0;bcd2<=2;bcd1<=8;bcd0<=4; end
			285: begin bcd3<=0;bcd2<=2;bcd1<=8;bcd0<=5; end
			286: begin bcd3<=0;bcd2<=2;bcd1<=8;bcd0<=6; end
			287: begin bcd3<=0;bcd2<=2;bcd1<=8;bcd0<=7; end
			288: begin bcd3<=0;bcd2<=2;bcd1<=8;bcd0<=8; end
			289: begin bcd3<=0;bcd2<=2;bcd1<=8;bcd0<=9; end
			290: begin bcd3<=0;bcd2<=2;bcd1<=9;bcd0<=0; end
			291: begin bcd3<=0;bcd2<=2;bcd1<=9;bcd0<=1; end
			292: begin bcd3<=0;bcd2<=2;bcd1<=9;bcd0<=2; end
			293: begin bcd3<=0;bcd2<=2;bcd1<=9;bcd0<=3; end
			294: begin bcd3<=0;bcd2<=2;bcd1<=9;bcd0<=4; end
			295: begin bcd3<=0;bcd2<=2;bcd1<=9;bcd0<=5; end
			296: begin bcd3<=0;bcd2<=2;bcd1<=9;bcd0<=6; end
			297: begin bcd3<=0;bcd2<=2;bcd1<=9;bcd0<=7; end
			298: begin bcd3<=0;bcd2<=2;bcd1<=9;bcd0<=8; end
			299: begin bcd3<=0;bcd2<=2;bcd1<=9;bcd0<=9; end
			300: begin bcd3<=0;bcd2<=3;bcd1<=0;bcd0<=0; end
			301: begin bcd3<=0;bcd2<=3;bcd1<=0;bcd0<=1; end
			302: begin bcd3<=0;bcd2<=3;bcd1<=0;bcd0<=2; end
			303: begin bcd3<=0;bcd2<=3;bcd1<=0;bcd0<=3; end
			304: begin bcd3<=0;bcd2<=3;bcd1<=0;bcd0<=4; end
			305: begin bcd3<=0;bcd2<=3;bcd1<=0;bcd0<=5; end
			306: begin bcd3<=0;bcd2<=3;bcd1<=0;bcd0<=6; end
			307: begin bcd3<=0;bcd2<=3;bcd1<=0;bcd0<=7; end
			308: begin bcd3<=0;bcd2<=3;bcd1<=0;bcd0<=8; end
			309: begin bcd3<=0;bcd2<=3;bcd1<=0;bcd0<=9; end
			310: begin bcd3<=0;bcd2<=3;bcd1<=1;bcd0<=0; end
			311: begin bcd3<=0;bcd2<=3;bcd1<=1;bcd0<=1; end
			312: begin bcd3<=0;bcd2<=3;bcd1<=1;bcd0<=2; end
			313: begin bcd3<=0;bcd2<=3;bcd1<=1;bcd0<=3; end
			314: begin bcd3<=0;bcd2<=3;bcd1<=1;bcd0<=4; end
			315: begin bcd3<=0;bcd2<=3;bcd1<=1;bcd0<=5; end
			316: begin bcd3<=0;bcd2<=3;bcd1<=1;bcd0<=6; end
			317: begin bcd3<=0;bcd2<=3;bcd1<=1;bcd0<=7; end
			318: begin bcd3<=0;bcd2<=3;bcd1<=1;bcd0<=8; end
			319: begin bcd3<=0;bcd2<=3;bcd1<=1;bcd0<=9; end
			320: begin bcd3<=0;bcd2<=3;bcd1<=2;bcd0<=0; end
			321: begin bcd3<=0;bcd2<=3;bcd1<=2;bcd0<=1; end
			322: begin bcd3<=0;bcd2<=3;bcd1<=2;bcd0<=2; end
			323: begin bcd3<=0;bcd2<=3;bcd1<=2;bcd0<=3; end
			324: begin bcd3<=0;bcd2<=3;bcd1<=2;bcd0<=4; end
			325: begin bcd3<=0;bcd2<=3;bcd1<=2;bcd0<=5; end
			326: begin bcd3<=0;bcd2<=3;bcd1<=2;bcd0<=6; end
			327: begin bcd3<=0;bcd2<=3;bcd1<=2;bcd0<=7; end
			328: begin bcd3<=0;bcd2<=3;bcd1<=2;bcd0<=8; end
			329: begin bcd3<=0;bcd2<=3;bcd1<=2;bcd0<=9; end
			330: begin bcd3<=0;bcd2<=3;bcd1<=3;bcd0<=0; end
			331: begin bcd3<=0;bcd2<=3;bcd1<=3;bcd0<=1; end
			332: begin bcd3<=0;bcd2<=3;bcd1<=3;bcd0<=2; end
			333: begin bcd3<=0;bcd2<=3;bcd1<=3;bcd0<=3; end
			334: begin bcd3<=0;bcd2<=3;bcd1<=3;bcd0<=4; end
			335: begin bcd3<=0;bcd2<=3;bcd1<=3;bcd0<=5; end
			336: begin bcd3<=0;bcd2<=3;bcd1<=3;bcd0<=6; end
			337: begin bcd3<=0;bcd2<=3;bcd1<=3;bcd0<=7; end
			338: begin bcd3<=0;bcd2<=3;bcd1<=3;bcd0<=8; end
			339: begin bcd3<=0;bcd2<=3;bcd1<=3;bcd0<=9; end
			340: begin bcd3<=0;bcd2<=3;bcd1<=4;bcd0<=0; end
			341: begin bcd3<=0;bcd2<=3;bcd1<=4;bcd0<=1; end
			342: begin bcd3<=0;bcd2<=3;bcd1<=4;bcd0<=2; end
			343: begin bcd3<=0;bcd2<=3;bcd1<=4;bcd0<=3; end
			344: begin bcd3<=0;bcd2<=3;bcd1<=4;bcd0<=4; end
			345: begin bcd3<=0;bcd2<=3;bcd1<=4;bcd0<=5; end
			346: begin bcd3<=0;bcd2<=3;bcd1<=4;bcd0<=6; end
			347: begin bcd3<=0;bcd2<=3;bcd1<=4;bcd0<=7; end
			348: begin bcd3<=0;bcd2<=3;bcd1<=4;bcd0<=8; end
			349: begin bcd3<=0;bcd2<=3;bcd1<=4;bcd0<=9; end
			350: begin bcd3<=0;bcd2<=3;bcd1<=5;bcd0<=0; end
			351: begin bcd3<=0;bcd2<=3;bcd1<=5;bcd0<=1; end
			352: begin bcd3<=0;bcd2<=3;bcd1<=5;bcd0<=2; end
			353: begin bcd3<=0;bcd2<=3;bcd1<=5;bcd0<=3; end
			354: begin bcd3<=0;bcd2<=3;bcd1<=5;bcd0<=4; end
			355: begin bcd3<=0;bcd2<=3;bcd1<=5;bcd0<=5; end
			356: begin bcd3<=0;bcd2<=3;bcd1<=5;bcd0<=6; end
			357: begin bcd3<=0;bcd2<=3;bcd1<=5;bcd0<=7; end
			358: begin bcd3<=0;bcd2<=3;bcd1<=5;bcd0<=8; end
			359: begin bcd3<=0;bcd2<=3;bcd1<=5;bcd0<=9; end
			360: begin bcd3<=0;bcd2<=3;bcd1<=6;bcd0<=0; end
			361: begin bcd3<=0;bcd2<=3;bcd1<=6;bcd0<=1; end
			362: begin bcd3<=0;bcd2<=3;bcd1<=6;bcd0<=2; end
			363: begin bcd3<=0;bcd2<=3;bcd1<=6;bcd0<=3; end
			364: begin bcd3<=0;bcd2<=3;bcd1<=6;bcd0<=4; end
			365: begin bcd3<=0;bcd2<=3;bcd1<=6;bcd0<=5; end
			366: begin bcd3<=0;bcd2<=3;bcd1<=6;bcd0<=6; end
			367: begin bcd3<=0;bcd2<=3;bcd1<=6;bcd0<=7; end
			368: begin bcd3<=0;bcd2<=3;bcd1<=6;bcd0<=8; end
			369: begin bcd3<=0;bcd2<=3;bcd1<=6;bcd0<=9; end
			370: begin bcd3<=0;bcd2<=3;bcd1<=7;bcd0<=0; end
			371: begin bcd3<=0;bcd2<=3;bcd1<=7;bcd0<=1; end
			372: begin bcd3<=0;bcd2<=3;bcd1<=7;bcd0<=2; end
			373: begin bcd3<=0;bcd2<=3;bcd1<=7;bcd0<=3; end
			374: begin bcd3<=0;bcd2<=3;bcd1<=7;bcd0<=4; end
			375: begin bcd3<=0;bcd2<=3;bcd1<=7;bcd0<=5; end
			376: begin bcd3<=0;bcd2<=3;bcd1<=7;bcd0<=6; end
			377: begin bcd3<=0;bcd2<=3;bcd1<=7;bcd0<=7; end
			378: begin bcd3<=0;bcd2<=3;bcd1<=7;bcd0<=8; end
			379: begin bcd3<=0;bcd2<=3;bcd1<=7;bcd0<=9; end
			380: begin bcd3<=0;bcd2<=3;bcd1<=8;bcd0<=0; end
			381: begin bcd3<=0;bcd2<=3;bcd1<=8;bcd0<=1; end
			382: begin bcd3<=0;bcd2<=3;bcd1<=8;bcd0<=2; end
			383: begin bcd3<=0;bcd2<=3;bcd1<=8;bcd0<=3; end
			384: begin bcd3<=0;bcd2<=3;bcd1<=8;bcd0<=4; end
			385: begin bcd3<=0;bcd2<=3;bcd1<=8;bcd0<=5; end
			386: begin bcd3<=0;bcd2<=3;bcd1<=8;bcd0<=6; end
			387: begin bcd3<=0;bcd2<=3;bcd1<=8;bcd0<=7; end
			388: begin bcd3<=0;bcd2<=3;bcd1<=8;bcd0<=8; end
			389: begin bcd3<=0;bcd2<=3;bcd1<=8;bcd0<=9; end
			390: begin bcd3<=0;bcd2<=3;bcd1<=9;bcd0<=0; end
			391: begin bcd3<=0;bcd2<=3;bcd1<=9;bcd0<=1; end
			392: begin bcd3<=0;bcd2<=3;bcd1<=9;bcd0<=2; end
			393: begin bcd3<=0;bcd2<=3;bcd1<=9;bcd0<=3; end
			394: begin bcd3<=0;bcd2<=3;bcd1<=9;bcd0<=4; end
			395: begin bcd3<=0;bcd2<=3;bcd1<=9;bcd0<=5; end
			396: begin bcd3<=0;bcd2<=3;bcd1<=9;bcd0<=6; end
			397: begin bcd3<=0;bcd2<=3;bcd1<=9;bcd0<=7; end
			398: begin bcd3<=0;bcd2<=3;bcd1<=9;bcd0<=8; end
			399: begin bcd3<=0;bcd2<=3;bcd1<=9;bcd0<=9; end
			400: begin bcd3<=0;bcd2<=4;bcd1<=0;bcd0<=0; end
			401: begin bcd3<=0;bcd2<=4;bcd1<=0;bcd0<=1; end
			402: begin bcd3<=0;bcd2<=4;bcd1<=0;bcd0<=2; end
			403: begin bcd3<=0;bcd2<=4;bcd1<=0;bcd0<=3; end
			404: begin bcd3<=0;bcd2<=4;bcd1<=0;bcd0<=4; end
			405: begin bcd3<=0;bcd2<=4;bcd1<=0;bcd0<=5; end
			406: begin bcd3<=0;bcd2<=4;bcd1<=0;bcd0<=6; end
			407: begin bcd3<=0;bcd2<=4;bcd1<=0;bcd0<=7; end
			408: begin bcd3<=0;bcd2<=4;bcd1<=0;bcd0<=8; end
			409: begin bcd3<=0;bcd2<=4;bcd1<=0;bcd0<=9; end
			410: begin bcd3<=0;bcd2<=4;bcd1<=1;bcd0<=0; end
			411: begin bcd3<=0;bcd2<=4;bcd1<=1;bcd0<=1; end
			412: begin bcd3<=0;bcd2<=4;bcd1<=1;bcd0<=2; end
			413: begin bcd3<=0;bcd2<=4;bcd1<=1;bcd0<=3; end
			414: begin bcd3<=0;bcd2<=4;bcd1<=1;bcd0<=4; end
			415: begin bcd3<=0;bcd2<=4;bcd1<=1;bcd0<=5; end
			416: begin bcd3<=0;bcd2<=4;bcd1<=1;bcd0<=6; end
			417: begin bcd3<=0;bcd2<=4;bcd1<=1;bcd0<=7; end
			418: begin bcd3<=0;bcd2<=4;bcd1<=1;bcd0<=8; end
			419: begin bcd3<=0;bcd2<=4;bcd1<=1;bcd0<=9; end
			420: begin bcd3<=0;bcd2<=4;bcd1<=2;bcd0<=0; end
			421: begin bcd3<=0;bcd2<=4;bcd1<=2;bcd0<=1; end
			422: begin bcd3<=0;bcd2<=4;bcd1<=2;bcd0<=2; end
			423: begin bcd3<=0;bcd2<=4;bcd1<=2;bcd0<=3; end
			424: begin bcd3<=0;bcd2<=4;bcd1<=2;bcd0<=4; end
			425: begin bcd3<=0;bcd2<=4;bcd1<=2;bcd0<=5; end
			426: begin bcd3<=0;bcd2<=4;bcd1<=2;bcd0<=6; end
			427: begin bcd3<=0;bcd2<=4;bcd1<=2;bcd0<=7; end
			428: begin bcd3<=0;bcd2<=4;bcd1<=2;bcd0<=8; end
			429: begin bcd3<=0;bcd2<=4;bcd1<=2;bcd0<=9; end
			430: begin bcd3<=0;bcd2<=4;bcd1<=3;bcd0<=0; end
			431: begin bcd3<=0;bcd2<=4;bcd1<=3;bcd0<=1; end
			432: begin bcd3<=0;bcd2<=4;bcd1<=3;bcd0<=2; end
			433: begin bcd3<=0;bcd2<=4;bcd1<=3;bcd0<=3; end
			434: begin bcd3<=0;bcd2<=4;bcd1<=3;bcd0<=4; end
			435: begin bcd3<=0;bcd2<=4;bcd1<=3;bcd0<=5; end
			436: begin bcd3<=0;bcd2<=4;bcd1<=3;bcd0<=6; end
			437: begin bcd3<=0;bcd2<=4;bcd1<=3;bcd0<=7; end
			438: begin bcd3<=0;bcd2<=4;bcd1<=3;bcd0<=8; end
			439: begin bcd3<=0;bcd2<=4;bcd1<=3;bcd0<=9; end
			440: begin bcd3<=0;bcd2<=4;bcd1<=4;bcd0<=0; end
			441: begin bcd3<=0;bcd2<=4;bcd1<=4;bcd0<=1; end
			442: begin bcd3<=0;bcd2<=4;bcd1<=4;bcd0<=2; end
			443: begin bcd3<=0;bcd2<=4;bcd1<=4;bcd0<=3; end
			444: begin bcd3<=0;bcd2<=4;bcd1<=4;bcd0<=4; end
			445: begin bcd3<=0;bcd2<=4;bcd1<=4;bcd0<=5; end
			446: begin bcd3<=0;bcd2<=4;bcd1<=4;bcd0<=6; end
			447: begin bcd3<=0;bcd2<=4;bcd1<=4;bcd0<=7; end
			448: begin bcd3<=0;bcd2<=4;bcd1<=4;bcd0<=8; end
			449: begin bcd3<=0;bcd2<=4;bcd1<=4;bcd0<=9; end
			450: begin bcd3<=0;bcd2<=4;bcd1<=5;bcd0<=0; end
			451: begin bcd3<=0;bcd2<=4;bcd1<=5;bcd0<=1; end
			452: begin bcd3<=0;bcd2<=4;bcd1<=5;bcd0<=2; end
			453: begin bcd3<=0;bcd2<=4;bcd1<=5;bcd0<=3; end
			454: begin bcd3<=0;bcd2<=4;bcd1<=5;bcd0<=4; end
			455: begin bcd3<=0;bcd2<=4;bcd1<=5;bcd0<=5; end
			456: begin bcd3<=0;bcd2<=4;bcd1<=5;bcd0<=6; end
			457: begin bcd3<=0;bcd2<=4;bcd1<=5;bcd0<=7; end
			458: begin bcd3<=0;bcd2<=4;bcd1<=5;bcd0<=8; end
			459: begin bcd3<=0;bcd2<=4;bcd1<=5;bcd0<=9; end
			460: begin bcd3<=0;bcd2<=4;bcd1<=6;bcd0<=0; end
			461: begin bcd3<=0;bcd2<=4;bcd1<=6;bcd0<=1; end
			462: begin bcd3<=0;bcd2<=4;bcd1<=6;bcd0<=2; end
			463: begin bcd3<=0;bcd2<=4;bcd1<=6;bcd0<=3; end
			464: begin bcd3<=0;bcd2<=4;bcd1<=6;bcd0<=4; end
			465: begin bcd3<=0;bcd2<=4;bcd1<=6;bcd0<=5; end
			466: begin bcd3<=0;bcd2<=4;bcd1<=6;bcd0<=6; end
			467: begin bcd3<=0;bcd2<=4;bcd1<=6;bcd0<=7; end
			468: begin bcd3<=0;bcd2<=4;bcd1<=6;bcd0<=8; end
			469: begin bcd3<=0;bcd2<=4;bcd1<=6;bcd0<=9; end
			470: begin bcd3<=0;bcd2<=4;bcd1<=7;bcd0<=0; end
			471: begin bcd3<=0;bcd2<=4;bcd1<=7;bcd0<=1; end
			472: begin bcd3<=0;bcd2<=4;bcd1<=7;bcd0<=2; end
			473: begin bcd3<=0;bcd2<=4;bcd1<=7;bcd0<=3; end
			474: begin bcd3<=0;bcd2<=4;bcd1<=7;bcd0<=4; end
			475: begin bcd3<=0;bcd2<=4;bcd1<=7;bcd0<=5; end
			476: begin bcd3<=0;bcd2<=4;bcd1<=7;bcd0<=6; end
			477: begin bcd3<=0;bcd2<=4;bcd1<=7;bcd0<=7; end
			478: begin bcd3<=0;bcd2<=4;bcd1<=7;bcd0<=8; end
			479: begin bcd3<=0;bcd2<=4;bcd1<=7;bcd0<=9; end
			480: begin bcd3<=0;bcd2<=4;bcd1<=8;bcd0<=0; end
			481: begin bcd3<=0;bcd2<=4;bcd1<=8;bcd0<=1; end
			482: begin bcd3<=0;bcd2<=4;bcd1<=8;bcd0<=2; end
			483: begin bcd3<=0;bcd2<=4;bcd1<=8;bcd0<=3; end
			484: begin bcd3<=0;bcd2<=4;bcd1<=8;bcd0<=4; end
			485: begin bcd3<=0;bcd2<=4;bcd1<=8;bcd0<=5; end
			486: begin bcd3<=0;bcd2<=4;bcd1<=8;bcd0<=6; end
			487: begin bcd3<=0;bcd2<=4;bcd1<=8;bcd0<=7; end
			488: begin bcd3<=0;bcd2<=4;bcd1<=8;bcd0<=8; end
			489: begin bcd3<=0;bcd2<=4;bcd1<=8;bcd0<=9; end
			490: begin bcd3<=0;bcd2<=4;bcd1<=9;bcd0<=0; end
			491: begin bcd3<=0;bcd2<=4;bcd1<=9;bcd0<=1; end
			492: begin bcd3<=0;bcd2<=4;bcd1<=9;bcd0<=2; end
			493: begin bcd3<=0;bcd2<=4;bcd1<=9;bcd0<=3; end
			494: begin bcd3<=0;bcd2<=4;bcd1<=9;bcd0<=4; end
			495: begin bcd3<=0;bcd2<=4;bcd1<=9;bcd0<=5; end
			496: begin bcd3<=0;bcd2<=4;bcd1<=9;bcd0<=6; end
			497: begin bcd3<=0;bcd2<=4;bcd1<=9;bcd0<=7; end
			498: begin bcd3<=0;bcd2<=4;bcd1<=9;bcd0<=8; end
			499: begin bcd3<=0;bcd2<=4;bcd1<=9;bcd0<=9; end
			500: begin bcd3<=0;bcd2<=5;bcd1<=0;bcd0<=0; end
			501: begin bcd3<=0;bcd2<=5;bcd1<=0;bcd0<=1; end
			502: begin bcd3<=0;bcd2<=5;bcd1<=0;bcd0<=2; end
			503: begin bcd3<=0;bcd2<=5;bcd1<=0;bcd0<=3; end
			504: begin bcd3<=0;bcd2<=5;bcd1<=0;bcd0<=4; end
			505: begin bcd3<=0;bcd2<=5;bcd1<=0;bcd0<=5; end
			506: begin bcd3<=0;bcd2<=5;bcd1<=0;bcd0<=6; end
			507: begin bcd3<=0;bcd2<=5;bcd1<=0;bcd0<=7; end
			508: begin bcd3<=0;bcd2<=5;bcd1<=0;bcd0<=8; end
			509: begin bcd3<=0;bcd2<=5;bcd1<=0;bcd0<=9; end
			510: begin bcd3<=0;bcd2<=5;bcd1<=1;bcd0<=0; end
			511: begin bcd3<=0;bcd2<=5;bcd1<=1;bcd0<=1; end
			512: begin bcd3<=0;bcd2<=5;bcd1<=1;bcd0<=2; end
			513: begin bcd3<=0;bcd2<=5;bcd1<=1;bcd0<=3; end
			514: begin bcd3<=0;bcd2<=5;bcd1<=1;bcd0<=4; end
			515: begin bcd3<=0;bcd2<=5;bcd1<=1;bcd0<=5; end
			516: begin bcd3<=0;bcd2<=5;bcd1<=1;bcd0<=6; end
			517: begin bcd3<=0;bcd2<=5;bcd1<=1;bcd0<=7; end
			518: begin bcd3<=0;bcd2<=5;bcd1<=1;bcd0<=8; end
			519: begin bcd3<=0;bcd2<=5;bcd1<=1;bcd0<=9; end
			520: begin bcd3<=0;bcd2<=5;bcd1<=2;bcd0<=0; end
			521: begin bcd3<=0;bcd2<=5;bcd1<=2;bcd0<=1; end
			522: begin bcd3<=0;bcd2<=5;bcd1<=2;bcd0<=2; end
			523: begin bcd3<=0;bcd2<=5;bcd1<=2;bcd0<=3; end
			524: begin bcd3<=0;bcd2<=5;bcd1<=2;bcd0<=4; end
			525: begin bcd3<=0;bcd2<=5;bcd1<=2;bcd0<=5; end
			526: begin bcd3<=0;bcd2<=5;bcd1<=2;bcd0<=6; end
			527: begin bcd3<=0;bcd2<=5;bcd1<=2;bcd0<=7; end
			528: begin bcd3<=0;bcd2<=5;bcd1<=2;bcd0<=8; end
			529: begin bcd3<=0;bcd2<=5;bcd1<=2;bcd0<=9; end
			530: begin bcd3<=0;bcd2<=5;bcd1<=3;bcd0<=0; end
			531: begin bcd3<=0;bcd2<=5;bcd1<=3;bcd0<=1; end
			532: begin bcd3<=0;bcd2<=5;bcd1<=3;bcd0<=2; end
			533: begin bcd3<=0;bcd2<=5;bcd1<=3;bcd0<=3; end
			534: begin bcd3<=0;bcd2<=5;bcd1<=3;bcd0<=4; end
			535: begin bcd3<=0;bcd2<=5;bcd1<=3;bcd0<=5; end
			536: begin bcd3<=0;bcd2<=5;bcd1<=3;bcd0<=6; end
			537: begin bcd3<=0;bcd2<=5;bcd1<=3;bcd0<=7; end
			538: begin bcd3<=0;bcd2<=5;bcd1<=3;bcd0<=8; end
			539: begin bcd3<=0;bcd2<=5;bcd1<=3;bcd0<=9; end
			540: begin bcd3<=0;bcd2<=5;bcd1<=4;bcd0<=0; end
			541: begin bcd3<=0;bcd2<=5;bcd1<=4;bcd0<=1; end
			542: begin bcd3<=0;bcd2<=5;bcd1<=4;bcd0<=2; end
			543: begin bcd3<=0;bcd2<=5;bcd1<=4;bcd0<=3; end
			544: begin bcd3<=0;bcd2<=5;bcd1<=4;bcd0<=4; end
			545: begin bcd3<=0;bcd2<=5;bcd1<=4;bcd0<=5; end
			546: begin bcd3<=0;bcd2<=5;bcd1<=4;bcd0<=6; end
			547: begin bcd3<=0;bcd2<=5;bcd1<=4;bcd0<=7; end
			548: begin bcd3<=0;bcd2<=5;bcd1<=4;bcd0<=8; end
			549: begin bcd3<=0;bcd2<=5;bcd1<=4;bcd0<=9; end
			550: begin bcd3<=0;bcd2<=5;bcd1<=5;bcd0<=0; end
			551: begin bcd3<=0;bcd2<=5;bcd1<=5;bcd0<=1; end
			552: begin bcd3<=0;bcd2<=5;bcd1<=5;bcd0<=2; end
			553: begin bcd3<=0;bcd2<=5;bcd1<=5;bcd0<=3; end
			554: begin bcd3<=0;bcd2<=5;bcd1<=5;bcd0<=4; end
			555: begin bcd3<=0;bcd2<=5;bcd1<=5;bcd0<=5; end
			556: begin bcd3<=0;bcd2<=5;bcd1<=5;bcd0<=6; end
			557: begin bcd3<=0;bcd2<=5;bcd1<=5;bcd0<=7; end
			558: begin bcd3<=0;bcd2<=5;bcd1<=5;bcd0<=8; end
			559: begin bcd3<=0;bcd2<=5;bcd1<=5;bcd0<=9; end
			560: begin bcd3<=0;bcd2<=5;bcd1<=6;bcd0<=0; end
			561: begin bcd3<=0;bcd2<=5;bcd1<=6;bcd0<=1; end
			562: begin bcd3<=0;bcd2<=5;bcd1<=6;bcd0<=2; end
			563: begin bcd3<=0;bcd2<=5;bcd1<=6;bcd0<=3; end
			564: begin bcd3<=0;bcd2<=5;bcd1<=6;bcd0<=4; end
			565: begin bcd3<=0;bcd2<=5;bcd1<=6;bcd0<=5; end
			566: begin bcd3<=0;bcd2<=5;bcd1<=6;bcd0<=6; end
			567: begin bcd3<=0;bcd2<=5;bcd1<=6;bcd0<=7; end
			568: begin bcd3<=0;bcd2<=5;bcd1<=6;bcd0<=8; end
			569: begin bcd3<=0;bcd2<=5;bcd1<=6;bcd0<=9; end
			570: begin bcd3<=0;bcd2<=5;bcd1<=7;bcd0<=0; end
			571: begin bcd3<=0;bcd2<=5;bcd1<=7;bcd0<=1; end
			572: begin bcd3<=0;bcd2<=5;bcd1<=7;bcd0<=2; end
			573: begin bcd3<=0;bcd2<=5;bcd1<=7;bcd0<=3; end
			574: begin bcd3<=0;bcd2<=5;bcd1<=7;bcd0<=4; end
			575: begin bcd3<=0;bcd2<=5;bcd1<=7;bcd0<=5; end
			576: begin bcd3<=0;bcd2<=5;bcd1<=7;bcd0<=6; end
			577: begin bcd3<=0;bcd2<=5;bcd1<=7;bcd0<=7; end
			578: begin bcd3<=0;bcd2<=5;bcd1<=7;bcd0<=8; end
			579: begin bcd3<=0;bcd2<=5;bcd1<=7;bcd0<=9; end
			580: begin bcd3<=0;bcd2<=5;bcd1<=8;bcd0<=0; end
			581: begin bcd3<=0;bcd2<=5;bcd1<=8;bcd0<=1; end
			582: begin bcd3<=0;bcd2<=5;bcd1<=8;bcd0<=2; end
			583: begin bcd3<=0;bcd2<=5;bcd1<=8;bcd0<=3; end
			584: begin bcd3<=0;bcd2<=5;bcd1<=8;bcd0<=4; end
			585: begin bcd3<=0;bcd2<=5;bcd1<=8;bcd0<=5; end
			586: begin bcd3<=0;bcd2<=5;bcd1<=8;bcd0<=6; end
			587: begin bcd3<=0;bcd2<=5;bcd1<=8;bcd0<=7; end
			588: begin bcd3<=0;bcd2<=5;bcd1<=8;bcd0<=8; end
			589: begin bcd3<=0;bcd2<=5;bcd1<=8;bcd0<=9; end
			590: begin bcd3<=0;bcd2<=5;bcd1<=9;bcd0<=0; end
			591: begin bcd3<=0;bcd2<=5;bcd1<=9;bcd0<=1; end
			592: begin bcd3<=0;bcd2<=5;bcd1<=9;bcd0<=2; end
			593: begin bcd3<=0;bcd2<=5;bcd1<=9;bcd0<=3; end
			594: begin bcd3<=0;bcd2<=5;bcd1<=9;bcd0<=4; end
			595: begin bcd3<=0;bcd2<=5;bcd1<=9;bcd0<=5; end
			596: begin bcd3<=0;bcd2<=5;bcd1<=9;bcd0<=6; end
			597: begin bcd3<=0;bcd2<=5;bcd1<=9;bcd0<=7; end
			598: begin bcd3<=0;bcd2<=5;bcd1<=9;bcd0<=8; end
			599: begin bcd3<=0;bcd2<=5;bcd1<=9;bcd0<=9; end
			600: begin bcd3<=0;bcd2<=6;bcd1<=0;bcd0<=0; end
			601: begin bcd3<=0;bcd2<=6;bcd1<=0;bcd0<=1; end
			602: begin bcd3<=0;bcd2<=6;bcd1<=0;bcd0<=2; end
			603: begin bcd3<=0;bcd2<=6;bcd1<=0;bcd0<=3; end
			604: begin bcd3<=0;bcd2<=6;bcd1<=0;bcd0<=4; end
			605: begin bcd3<=0;bcd2<=6;bcd1<=0;bcd0<=5; end
			606: begin bcd3<=0;bcd2<=6;bcd1<=0;bcd0<=6; end
			607: begin bcd3<=0;bcd2<=6;bcd1<=0;bcd0<=7; end
			608: begin bcd3<=0;bcd2<=6;bcd1<=0;bcd0<=8; end
			609: begin bcd3<=0;bcd2<=6;bcd1<=0;bcd0<=9; end
			610: begin bcd3<=0;bcd2<=6;bcd1<=1;bcd0<=0; end
			611: begin bcd3<=0;bcd2<=6;bcd1<=1;bcd0<=1; end
			612: begin bcd3<=0;bcd2<=6;bcd1<=1;bcd0<=2; end
			613: begin bcd3<=0;bcd2<=6;bcd1<=1;bcd0<=3; end
			614: begin bcd3<=0;bcd2<=6;bcd1<=1;bcd0<=4; end
			615: begin bcd3<=0;bcd2<=6;bcd1<=1;bcd0<=5; end
			616: begin bcd3<=0;bcd2<=6;bcd1<=1;bcd0<=6; end
			617: begin bcd3<=0;bcd2<=6;bcd1<=1;bcd0<=7; end
			618: begin bcd3<=0;bcd2<=6;bcd1<=1;bcd0<=8; end
			619: begin bcd3<=0;bcd2<=6;bcd1<=1;bcd0<=9; end
			620: begin bcd3<=0;bcd2<=6;bcd1<=2;bcd0<=0; end
			621: begin bcd3<=0;bcd2<=6;bcd1<=2;bcd0<=1; end
			622: begin bcd3<=0;bcd2<=6;bcd1<=2;bcd0<=2; end
			623: begin bcd3<=0;bcd2<=6;bcd1<=2;bcd0<=3; end
			624: begin bcd3<=0;bcd2<=6;bcd1<=2;bcd0<=4; end
			625: begin bcd3<=0;bcd2<=6;bcd1<=2;bcd0<=5; end
			626: begin bcd3<=0;bcd2<=6;bcd1<=2;bcd0<=6; end
			627: begin bcd3<=0;bcd2<=6;bcd1<=2;bcd0<=7; end
			628: begin bcd3<=0;bcd2<=6;bcd1<=2;bcd0<=8; end
			629: begin bcd3<=0;bcd2<=6;bcd1<=2;bcd0<=9; end
			630: begin bcd3<=0;bcd2<=6;bcd1<=3;bcd0<=0; end
			631: begin bcd3<=0;bcd2<=6;bcd1<=3;bcd0<=1; end
			632: begin bcd3<=0;bcd2<=6;bcd1<=3;bcd0<=2; end
			633: begin bcd3<=0;bcd2<=6;bcd1<=3;bcd0<=3; end
			634: begin bcd3<=0;bcd2<=6;bcd1<=3;bcd0<=4; end
			635: begin bcd3<=0;bcd2<=6;bcd1<=3;bcd0<=5; end
			636: begin bcd3<=0;bcd2<=6;bcd1<=3;bcd0<=6; end
			637: begin bcd3<=0;bcd2<=6;bcd1<=3;bcd0<=7; end
			638: begin bcd3<=0;bcd2<=6;bcd1<=3;bcd0<=8; end
			639: begin bcd3<=0;bcd2<=6;bcd1<=3;bcd0<=9; end
			640: begin bcd3<=0;bcd2<=6;bcd1<=4;bcd0<=0; end
			641: begin bcd3<=0;bcd2<=6;bcd1<=4;bcd0<=1; end
			642: begin bcd3<=0;bcd2<=6;bcd1<=4;bcd0<=2; end
			643: begin bcd3<=0;bcd2<=6;bcd1<=4;bcd0<=3; end
			644: begin bcd3<=0;bcd2<=6;bcd1<=4;bcd0<=4; end
			645: begin bcd3<=0;bcd2<=6;bcd1<=4;bcd0<=5; end
			646: begin bcd3<=0;bcd2<=6;bcd1<=4;bcd0<=6; end
			647: begin bcd3<=0;bcd2<=6;bcd1<=4;bcd0<=7; end
			648: begin bcd3<=0;bcd2<=6;bcd1<=4;bcd0<=8; end
			649: begin bcd3<=0;bcd2<=6;bcd1<=4;bcd0<=9; end
			650: begin bcd3<=0;bcd2<=6;bcd1<=5;bcd0<=0; end
			651: begin bcd3<=0;bcd2<=6;bcd1<=5;bcd0<=1; end
			652: begin bcd3<=0;bcd2<=6;bcd1<=5;bcd0<=2; end
			653: begin bcd3<=0;bcd2<=6;bcd1<=5;bcd0<=3; end
			654: begin bcd3<=0;bcd2<=6;bcd1<=5;bcd0<=4; end
			655: begin bcd3<=0;bcd2<=6;bcd1<=5;bcd0<=5; end
			656: begin bcd3<=0;bcd2<=6;bcd1<=5;bcd0<=6; end
			657: begin bcd3<=0;bcd2<=6;bcd1<=5;bcd0<=7; end
			658: begin bcd3<=0;bcd2<=6;bcd1<=5;bcd0<=8; end
			659: begin bcd3<=0;bcd2<=6;bcd1<=5;bcd0<=9; end
			660: begin bcd3<=0;bcd2<=6;bcd1<=6;bcd0<=0; end
			661: begin bcd3<=0;bcd2<=6;bcd1<=6;bcd0<=1; end
			662: begin bcd3<=0;bcd2<=6;bcd1<=6;bcd0<=2; end
			663: begin bcd3<=0;bcd2<=6;bcd1<=6;bcd0<=3; end
			664: begin bcd3<=0;bcd2<=6;bcd1<=6;bcd0<=4; end
			665: begin bcd3<=0;bcd2<=6;bcd1<=6;bcd0<=5; end
			666: begin bcd3<=0;bcd2<=6;bcd1<=6;bcd0<=6; end
			667: begin bcd3<=0;bcd2<=6;bcd1<=6;bcd0<=7; end
			668: begin bcd3<=0;bcd2<=6;bcd1<=6;bcd0<=8; end
			669: begin bcd3<=0;bcd2<=6;bcd1<=6;bcd0<=9; end
			670: begin bcd3<=0;bcd2<=6;bcd1<=7;bcd0<=0; end
			671: begin bcd3<=0;bcd2<=6;bcd1<=7;bcd0<=1; end
			672: begin bcd3<=0;bcd2<=6;bcd1<=7;bcd0<=2; end
			673: begin bcd3<=0;bcd2<=6;bcd1<=7;bcd0<=3; end
			674: begin bcd3<=0;bcd2<=6;bcd1<=7;bcd0<=4; end
			675: begin bcd3<=0;bcd2<=6;bcd1<=7;bcd0<=5; end
			676: begin bcd3<=0;bcd2<=6;bcd1<=7;bcd0<=6; end
			677: begin bcd3<=0;bcd2<=6;bcd1<=7;bcd0<=7; end
			678: begin bcd3<=0;bcd2<=6;bcd1<=7;bcd0<=8; end
			679: begin bcd3<=0;bcd2<=6;bcd1<=7;bcd0<=9; end
			680: begin bcd3<=0;bcd2<=6;bcd1<=8;bcd0<=0; end
			681: begin bcd3<=0;bcd2<=6;bcd1<=8;bcd0<=1; end
			682: begin bcd3<=0;bcd2<=6;bcd1<=8;bcd0<=2; end
			683: begin bcd3<=0;bcd2<=6;bcd1<=8;bcd0<=3; end
			684: begin bcd3<=0;bcd2<=6;bcd1<=8;bcd0<=4; end
			685: begin bcd3<=0;bcd2<=6;bcd1<=8;bcd0<=5; end
			686: begin bcd3<=0;bcd2<=6;bcd1<=8;bcd0<=6; end
			687: begin bcd3<=0;bcd2<=6;bcd1<=8;bcd0<=7; end
			688: begin bcd3<=0;bcd2<=6;bcd1<=8;bcd0<=8; end
			689: begin bcd3<=0;bcd2<=6;bcd1<=8;bcd0<=9; end
			690: begin bcd3<=0;bcd2<=6;bcd1<=9;bcd0<=0; end
			691: begin bcd3<=0;bcd2<=6;bcd1<=9;bcd0<=1; end
			692: begin bcd3<=0;bcd2<=6;bcd1<=9;bcd0<=2; end
			693: begin bcd3<=0;bcd2<=6;bcd1<=9;bcd0<=3; end
			694: begin bcd3<=0;bcd2<=6;bcd1<=9;bcd0<=4; end
			695: begin bcd3<=0;bcd2<=6;bcd1<=9;bcd0<=5; end
			696: begin bcd3<=0;bcd2<=6;bcd1<=9;bcd0<=6; end
			697: begin bcd3<=0;bcd2<=6;bcd1<=9;bcd0<=7; end
			698: begin bcd3<=0;bcd2<=6;bcd1<=9;bcd0<=8; end
			699: begin bcd3<=0;bcd2<=6;bcd1<=9;bcd0<=9; end
			700: begin bcd3<=0;bcd2<=7;bcd1<=0;bcd0<=0; end
			701: begin bcd3<=0;bcd2<=7;bcd1<=0;bcd0<=1; end
			702: begin bcd3<=0;bcd2<=7;bcd1<=0;bcd0<=2; end
			703: begin bcd3<=0;bcd2<=7;bcd1<=0;bcd0<=3; end
			704: begin bcd3<=0;bcd2<=7;bcd1<=0;bcd0<=4; end
			705: begin bcd3<=0;bcd2<=7;bcd1<=0;bcd0<=5; end
			706: begin bcd3<=0;bcd2<=7;bcd1<=0;bcd0<=6; end
			707: begin bcd3<=0;bcd2<=7;bcd1<=0;bcd0<=7; end
			708: begin bcd3<=0;bcd2<=7;bcd1<=0;bcd0<=8; end
			709: begin bcd3<=0;bcd2<=7;bcd1<=0;bcd0<=9; end
			710: begin bcd3<=0;bcd2<=7;bcd1<=1;bcd0<=0; end
			711: begin bcd3<=0;bcd2<=7;bcd1<=1;bcd0<=1; end
			712: begin bcd3<=0;bcd2<=7;bcd1<=1;bcd0<=2; end
			713: begin bcd3<=0;bcd2<=7;bcd1<=1;bcd0<=3; end
			714: begin bcd3<=0;bcd2<=7;bcd1<=1;bcd0<=4; end
			715: begin bcd3<=0;bcd2<=7;bcd1<=1;bcd0<=5; end
			716: begin bcd3<=0;bcd2<=7;bcd1<=1;bcd0<=6; end
			717: begin bcd3<=0;bcd2<=7;bcd1<=1;bcd0<=7; end
			718: begin bcd3<=0;bcd2<=7;bcd1<=1;bcd0<=8; end
			719: begin bcd3<=0;bcd2<=7;bcd1<=1;bcd0<=9; end
			720: begin bcd3<=0;bcd2<=7;bcd1<=2;bcd0<=0; end
			721: begin bcd3<=0;bcd2<=7;bcd1<=2;bcd0<=1; end
			722: begin bcd3<=0;bcd2<=7;bcd1<=2;bcd0<=2; end
			723: begin bcd3<=0;bcd2<=7;bcd1<=2;bcd0<=3; end
			724: begin bcd3<=0;bcd2<=7;bcd1<=2;bcd0<=4; end
			725: begin bcd3<=0;bcd2<=7;bcd1<=2;bcd0<=5; end
			726: begin bcd3<=0;bcd2<=7;bcd1<=2;bcd0<=6; end
			727: begin bcd3<=0;bcd2<=7;bcd1<=2;bcd0<=7; end
			728: begin bcd3<=0;bcd2<=7;bcd1<=2;bcd0<=8; end
			729: begin bcd3<=0;bcd2<=7;bcd1<=2;bcd0<=9; end
			730: begin bcd3<=0;bcd2<=7;bcd1<=3;bcd0<=0; end
			731: begin bcd3<=0;bcd2<=7;bcd1<=3;bcd0<=1; end
			732: begin bcd3<=0;bcd2<=7;bcd1<=3;bcd0<=2; end
			733: begin bcd3<=0;bcd2<=7;bcd1<=3;bcd0<=3; end
			734: begin bcd3<=0;bcd2<=7;bcd1<=3;bcd0<=4; end
			735: begin bcd3<=0;bcd2<=7;bcd1<=3;bcd0<=5; end
			736: begin bcd3<=0;bcd2<=7;bcd1<=3;bcd0<=6; end
			737: begin bcd3<=0;bcd2<=7;bcd1<=3;bcd0<=7; end
			738: begin bcd3<=0;bcd2<=7;bcd1<=3;bcd0<=8; end
			739: begin bcd3<=0;bcd2<=7;bcd1<=3;bcd0<=9; end
			740: begin bcd3<=0;bcd2<=7;bcd1<=4;bcd0<=0; end
			741: begin bcd3<=0;bcd2<=7;bcd1<=4;bcd0<=1; end
			742: begin bcd3<=0;bcd2<=7;bcd1<=4;bcd0<=2; end
			743: begin bcd3<=0;bcd2<=7;bcd1<=4;bcd0<=3; end
			744: begin bcd3<=0;bcd2<=7;bcd1<=4;bcd0<=4; end
			745: begin bcd3<=0;bcd2<=7;bcd1<=4;bcd0<=5; end
			746: begin bcd3<=0;bcd2<=7;bcd1<=4;bcd0<=6; end
			747: begin bcd3<=0;bcd2<=7;bcd1<=4;bcd0<=7; end
			748: begin bcd3<=0;bcd2<=7;bcd1<=4;bcd0<=8; end
			749: begin bcd3<=0;bcd2<=7;bcd1<=4;bcd0<=9; end
			750: begin bcd3<=0;bcd2<=7;bcd1<=5;bcd0<=0; end
			751: begin bcd3<=0;bcd2<=7;bcd1<=5;bcd0<=1; end
			752: begin bcd3<=0;bcd2<=7;bcd1<=5;bcd0<=2; end
			753: begin bcd3<=0;bcd2<=7;bcd1<=5;bcd0<=3; end
			754: begin bcd3<=0;bcd2<=7;bcd1<=5;bcd0<=4; end
			755: begin bcd3<=0;bcd2<=7;bcd1<=5;bcd0<=5; end
			756: begin bcd3<=0;bcd2<=7;bcd1<=5;bcd0<=6; end
			757: begin bcd3<=0;bcd2<=7;bcd1<=5;bcd0<=7; end
			758: begin bcd3<=0;bcd2<=7;bcd1<=5;bcd0<=8; end
			759: begin bcd3<=0;bcd2<=7;bcd1<=5;bcd0<=9; end
			760: begin bcd3<=0;bcd2<=7;bcd1<=6;bcd0<=0; end
			761: begin bcd3<=0;bcd2<=7;bcd1<=6;bcd0<=1; end
			762: begin bcd3<=0;bcd2<=7;bcd1<=6;bcd0<=2; end
			763: begin bcd3<=0;bcd2<=7;bcd1<=6;bcd0<=3; end
			764: begin bcd3<=0;bcd2<=7;bcd1<=6;bcd0<=4; end
			765: begin bcd3<=0;bcd2<=7;bcd1<=6;bcd0<=5; end
			766: begin bcd3<=0;bcd2<=7;bcd1<=6;bcd0<=6; end
			767: begin bcd3<=0;bcd2<=7;bcd1<=6;bcd0<=7; end
			768: begin bcd3<=0;bcd2<=7;bcd1<=6;bcd0<=8; end
			769: begin bcd3<=0;bcd2<=7;bcd1<=6;bcd0<=9; end
			770: begin bcd3<=0;bcd2<=7;bcd1<=7;bcd0<=0; end
			771: begin bcd3<=0;bcd2<=7;bcd1<=7;bcd0<=1; end
			772: begin bcd3<=0;bcd2<=7;bcd1<=7;bcd0<=2; end
			773: begin bcd3<=0;bcd2<=7;bcd1<=7;bcd0<=3; end
			774: begin bcd3<=0;bcd2<=7;bcd1<=7;bcd0<=4; end
			775: begin bcd3<=0;bcd2<=7;bcd1<=7;bcd0<=5; end
			776: begin bcd3<=0;bcd2<=7;bcd1<=7;bcd0<=6; end
			777: begin bcd3<=0;bcd2<=7;bcd1<=7;bcd0<=7; end
			778: begin bcd3<=0;bcd2<=7;bcd1<=7;bcd0<=8; end
			779: begin bcd3<=0;bcd2<=7;bcd1<=7;bcd0<=9; end
			780: begin bcd3<=0;bcd2<=7;bcd1<=8;bcd0<=0; end
			781: begin bcd3<=0;bcd2<=7;bcd1<=8;bcd0<=1; end
			782: begin bcd3<=0;bcd2<=7;bcd1<=8;bcd0<=2; end
			783: begin bcd3<=0;bcd2<=7;bcd1<=8;bcd0<=3; end
			784: begin bcd3<=0;bcd2<=7;bcd1<=8;bcd0<=4; end
			785: begin bcd3<=0;bcd2<=7;bcd1<=8;bcd0<=5; end
			786: begin bcd3<=0;bcd2<=7;bcd1<=8;bcd0<=6; end
			787: begin bcd3<=0;bcd2<=7;bcd1<=8;bcd0<=7; end
			788: begin bcd3<=0;bcd2<=7;bcd1<=8;bcd0<=8; end
			789: begin bcd3<=0;bcd2<=7;bcd1<=8;bcd0<=9; end
			790: begin bcd3<=0;bcd2<=7;bcd1<=9;bcd0<=0; end
			791: begin bcd3<=0;bcd2<=7;bcd1<=9;bcd0<=1; end
			792: begin bcd3<=0;bcd2<=7;bcd1<=9;bcd0<=2; end
			793: begin bcd3<=0;bcd2<=7;bcd1<=9;bcd0<=3; end
			794: begin bcd3<=0;bcd2<=7;bcd1<=9;bcd0<=4; end
			795: begin bcd3<=0;bcd2<=7;bcd1<=9;bcd0<=5; end
			796: begin bcd3<=0;bcd2<=7;bcd1<=9;bcd0<=6; end
			797: begin bcd3<=0;bcd2<=7;bcd1<=9;bcd0<=7; end
			798: begin bcd3<=0;bcd2<=7;bcd1<=9;bcd0<=8; end
			799: begin bcd3<=0;bcd2<=7;bcd1<=9;bcd0<=9; end
			800: begin bcd3<=0;bcd2<=8;bcd1<=0;bcd0<=0; end
			801: begin bcd3<=0;bcd2<=8;bcd1<=0;bcd0<=1; end
			802: begin bcd3<=0;bcd2<=8;bcd1<=0;bcd0<=2; end
			803: begin bcd3<=0;bcd2<=8;bcd1<=0;bcd0<=3; end
			804: begin bcd3<=0;bcd2<=8;bcd1<=0;bcd0<=4; end
			805: begin bcd3<=0;bcd2<=8;bcd1<=0;bcd0<=5; end
			806: begin bcd3<=0;bcd2<=8;bcd1<=0;bcd0<=6; end
			807: begin bcd3<=0;bcd2<=8;bcd1<=0;bcd0<=7; end
			808: begin bcd3<=0;bcd2<=8;bcd1<=0;bcd0<=8; end
			809: begin bcd3<=0;bcd2<=8;bcd1<=0;bcd0<=9; end
			810: begin bcd3<=0;bcd2<=8;bcd1<=1;bcd0<=0; end
			811: begin bcd3<=0;bcd2<=8;bcd1<=1;bcd0<=1; end
			812: begin bcd3<=0;bcd2<=8;bcd1<=1;bcd0<=2; end
			813: begin bcd3<=0;bcd2<=8;bcd1<=1;bcd0<=3; end
			814: begin bcd3<=0;bcd2<=8;bcd1<=1;bcd0<=4; end
			815: begin bcd3<=0;bcd2<=8;bcd1<=1;bcd0<=5; end
			816: begin bcd3<=0;bcd2<=8;bcd1<=1;bcd0<=6; end
			817: begin bcd3<=0;bcd2<=8;bcd1<=1;bcd0<=7; end
			818: begin bcd3<=0;bcd2<=8;bcd1<=1;bcd0<=8; end
			819: begin bcd3<=0;bcd2<=8;bcd1<=1;bcd0<=9; end
			820: begin bcd3<=0;bcd2<=8;bcd1<=2;bcd0<=0; end
			821: begin bcd3<=0;bcd2<=8;bcd1<=2;bcd0<=1; end
			822: begin bcd3<=0;bcd2<=8;bcd1<=2;bcd0<=2; end
			823: begin bcd3<=0;bcd2<=8;bcd1<=2;bcd0<=3; end
			824: begin bcd3<=0;bcd2<=8;bcd1<=2;bcd0<=4; end
			825: begin bcd3<=0;bcd2<=8;bcd1<=2;bcd0<=5; end
			826: begin bcd3<=0;bcd2<=8;bcd1<=2;bcd0<=6; end
			827: begin bcd3<=0;bcd2<=8;bcd1<=2;bcd0<=7; end
			828: begin bcd3<=0;bcd2<=8;bcd1<=2;bcd0<=8; end
			829: begin bcd3<=0;bcd2<=8;bcd1<=2;bcd0<=9; end
			830: begin bcd3<=0;bcd2<=8;bcd1<=3;bcd0<=0; end
			831: begin bcd3<=0;bcd2<=8;bcd1<=3;bcd0<=1; end
			832: begin bcd3<=0;bcd2<=8;bcd1<=3;bcd0<=2; end
			833: begin bcd3<=0;bcd2<=8;bcd1<=3;bcd0<=3; end
			834: begin bcd3<=0;bcd2<=8;bcd1<=3;bcd0<=4; end
			835: begin bcd3<=0;bcd2<=8;bcd1<=3;bcd0<=5; end
			836: begin bcd3<=0;bcd2<=8;bcd1<=3;bcd0<=6; end
			837: begin bcd3<=0;bcd2<=8;bcd1<=3;bcd0<=7; end
			838: begin bcd3<=0;bcd2<=8;bcd1<=3;bcd0<=8; end
			839: begin bcd3<=0;bcd2<=8;bcd1<=3;bcd0<=9; end
			840: begin bcd3<=0;bcd2<=8;bcd1<=4;bcd0<=0; end
			841: begin bcd3<=0;bcd2<=8;bcd1<=4;bcd0<=1; end
			842: begin bcd3<=0;bcd2<=8;bcd1<=4;bcd0<=2; end
			843: begin bcd3<=0;bcd2<=8;bcd1<=4;bcd0<=3; end
			844: begin bcd3<=0;bcd2<=8;bcd1<=4;bcd0<=4; end
			845: begin bcd3<=0;bcd2<=8;bcd1<=4;bcd0<=5; end
			846: begin bcd3<=0;bcd2<=8;bcd1<=4;bcd0<=6; end
			847: begin bcd3<=0;bcd2<=8;bcd1<=4;bcd0<=7; end
			848: begin bcd3<=0;bcd2<=8;bcd1<=4;bcd0<=8; end
			849: begin bcd3<=0;bcd2<=8;bcd1<=4;bcd0<=9; end
			850: begin bcd3<=0;bcd2<=8;bcd1<=5;bcd0<=0; end
			851: begin bcd3<=0;bcd2<=8;bcd1<=5;bcd0<=1; end
			852: begin bcd3<=0;bcd2<=8;bcd1<=5;bcd0<=2; end
			853: begin bcd3<=0;bcd2<=8;bcd1<=5;bcd0<=3; end
			854: begin bcd3<=0;bcd2<=8;bcd1<=5;bcd0<=4; end
			855: begin bcd3<=0;bcd2<=8;bcd1<=5;bcd0<=5; end
			856: begin bcd3<=0;bcd2<=8;bcd1<=5;bcd0<=6; end
			857: begin bcd3<=0;bcd2<=8;bcd1<=5;bcd0<=7; end
			858: begin bcd3<=0;bcd2<=8;bcd1<=5;bcd0<=8; end
			859: begin bcd3<=0;bcd2<=8;bcd1<=5;bcd0<=9; end
			860: begin bcd3<=0;bcd2<=8;bcd1<=6;bcd0<=0; end
			861: begin bcd3<=0;bcd2<=8;bcd1<=6;bcd0<=1; end
			862: begin bcd3<=0;bcd2<=8;bcd1<=6;bcd0<=2; end
			863: begin bcd3<=0;bcd2<=8;bcd1<=6;bcd0<=3; end
			864: begin bcd3<=0;bcd2<=8;bcd1<=6;bcd0<=4; end
			865: begin bcd3<=0;bcd2<=8;bcd1<=6;bcd0<=5; end
			866: begin bcd3<=0;bcd2<=8;bcd1<=6;bcd0<=6; end
			867: begin bcd3<=0;bcd2<=8;bcd1<=6;bcd0<=7; end
			868: begin bcd3<=0;bcd2<=8;bcd1<=6;bcd0<=8; end
			869: begin bcd3<=0;bcd2<=8;bcd1<=6;bcd0<=9; end
			870: begin bcd3<=0;bcd2<=8;bcd1<=7;bcd0<=0; end
			871: begin bcd3<=0;bcd2<=8;bcd1<=7;bcd0<=1; end
			872: begin bcd3<=0;bcd2<=8;bcd1<=7;bcd0<=2; end
			873: begin bcd3<=0;bcd2<=8;bcd1<=7;bcd0<=3; end
			874: begin bcd3<=0;bcd2<=8;bcd1<=7;bcd0<=4; end
			875: begin bcd3<=0;bcd2<=8;bcd1<=7;bcd0<=5; end
			876: begin bcd3<=0;bcd2<=8;bcd1<=7;bcd0<=6; end
			877: begin bcd3<=0;bcd2<=8;bcd1<=7;bcd0<=7; end
			878: begin bcd3<=0;bcd2<=8;bcd1<=7;bcd0<=8; end
			879: begin bcd3<=0;bcd2<=8;bcd1<=7;bcd0<=9; end
			880: begin bcd3<=0;bcd2<=8;bcd1<=8;bcd0<=0; end
			881: begin bcd3<=0;bcd2<=8;bcd1<=8;bcd0<=1; end
			882: begin bcd3<=0;bcd2<=8;bcd1<=8;bcd0<=2; end
			883: begin bcd3<=0;bcd2<=8;bcd1<=8;bcd0<=3; end
			884: begin bcd3<=0;bcd2<=8;bcd1<=8;bcd0<=4; end
			885: begin bcd3<=0;bcd2<=8;bcd1<=8;bcd0<=5; end
			886: begin bcd3<=0;bcd2<=8;bcd1<=8;bcd0<=6; end
			887: begin bcd3<=0;bcd2<=8;bcd1<=8;bcd0<=7; end
			888: begin bcd3<=0;bcd2<=8;bcd1<=8;bcd0<=8; end
			889: begin bcd3<=0;bcd2<=8;bcd1<=8;bcd0<=9; end
			890: begin bcd3<=0;bcd2<=8;bcd1<=9;bcd0<=0; end
			891: begin bcd3<=0;bcd2<=8;bcd1<=9;bcd0<=1; end
			892: begin bcd3<=0;bcd2<=8;bcd1<=9;bcd0<=2; end
			893: begin bcd3<=0;bcd2<=8;bcd1<=9;bcd0<=3; end
			894: begin bcd3<=0;bcd2<=8;bcd1<=9;bcd0<=4; end
			895: begin bcd3<=0;bcd2<=8;bcd1<=9;bcd0<=5; end
			896: begin bcd3<=0;bcd2<=8;bcd1<=9;bcd0<=6; end
			897: begin bcd3<=0;bcd2<=8;bcd1<=9;bcd0<=7; end
			898: begin bcd3<=0;bcd2<=8;bcd1<=9;bcd0<=8; end
			899: begin bcd3<=0;bcd2<=8;bcd1<=9;bcd0<=9; end
			900: begin bcd3<=0;bcd2<=9;bcd1<=0;bcd0<=0; end
			901: begin bcd3<=0;bcd2<=9;bcd1<=0;bcd0<=1; end
			902: begin bcd3<=0;bcd2<=9;bcd1<=0;bcd0<=2; end
			903: begin bcd3<=0;bcd2<=9;bcd1<=0;bcd0<=3; end
			904: begin bcd3<=0;bcd2<=9;bcd1<=0;bcd0<=4; end
			905: begin bcd3<=0;bcd2<=9;bcd1<=0;bcd0<=5; end
			906: begin bcd3<=0;bcd2<=9;bcd1<=0;bcd0<=6; end
			907: begin bcd3<=0;bcd2<=9;bcd1<=0;bcd0<=7; end
			908: begin bcd3<=0;bcd2<=9;bcd1<=0;bcd0<=8; end
			909: begin bcd3<=0;bcd2<=9;bcd1<=0;bcd0<=9; end
			910: begin bcd3<=0;bcd2<=9;bcd1<=1;bcd0<=0; end
			911: begin bcd3<=0;bcd2<=9;bcd1<=1;bcd0<=1; end
			912: begin bcd3<=0;bcd2<=9;bcd1<=1;bcd0<=2; end
			913: begin bcd3<=0;bcd2<=9;bcd1<=1;bcd0<=3; end
			914: begin bcd3<=0;bcd2<=9;bcd1<=1;bcd0<=4; end
			915: begin bcd3<=0;bcd2<=9;bcd1<=1;bcd0<=5; end
			916: begin bcd3<=0;bcd2<=9;bcd1<=1;bcd0<=6; end
			917: begin bcd3<=0;bcd2<=9;bcd1<=1;bcd0<=7; end
			918: begin bcd3<=0;bcd2<=9;bcd1<=1;bcd0<=8; end
			919: begin bcd3<=0;bcd2<=9;bcd1<=1;bcd0<=9; end
			920: begin bcd3<=0;bcd2<=9;bcd1<=2;bcd0<=0; end
			921: begin bcd3<=0;bcd2<=9;bcd1<=2;bcd0<=1; end
			922: begin bcd3<=0;bcd2<=9;bcd1<=2;bcd0<=2; end
			923: begin bcd3<=0;bcd2<=9;bcd1<=2;bcd0<=3; end
			924: begin bcd3<=0;bcd2<=9;bcd1<=2;bcd0<=4; end
			925: begin bcd3<=0;bcd2<=9;bcd1<=2;bcd0<=5; end
			926: begin bcd3<=0;bcd2<=9;bcd1<=2;bcd0<=6; end
			927: begin bcd3<=0;bcd2<=9;bcd1<=2;bcd0<=7; end
			928: begin bcd3<=0;bcd2<=9;bcd1<=2;bcd0<=8; end
			929: begin bcd3<=0;bcd2<=9;bcd1<=2;bcd0<=9; end
			930: begin bcd3<=0;bcd2<=9;bcd1<=3;bcd0<=0; end
			931: begin bcd3<=0;bcd2<=9;bcd1<=3;bcd0<=1; end
			932: begin bcd3<=0;bcd2<=9;bcd1<=3;bcd0<=2; end
			933: begin bcd3<=0;bcd2<=9;bcd1<=3;bcd0<=3; end
			934: begin bcd3<=0;bcd2<=9;bcd1<=3;bcd0<=4; end
			935: begin bcd3<=0;bcd2<=9;bcd1<=3;bcd0<=5; end
			936: begin bcd3<=0;bcd2<=9;bcd1<=3;bcd0<=6; end
			937: begin bcd3<=0;bcd2<=9;bcd1<=3;bcd0<=7; end
			938: begin bcd3<=0;bcd2<=9;bcd1<=3;bcd0<=8; end
			939: begin bcd3<=0;bcd2<=9;bcd1<=3;bcd0<=9; end
			940: begin bcd3<=0;bcd2<=9;bcd1<=4;bcd0<=0; end
			941: begin bcd3<=0;bcd2<=9;bcd1<=4;bcd0<=1; end
			942: begin bcd3<=0;bcd2<=9;bcd1<=4;bcd0<=2; end
			943: begin bcd3<=0;bcd2<=9;bcd1<=4;bcd0<=3; end
			944: begin bcd3<=0;bcd2<=9;bcd1<=4;bcd0<=4; end
			945: begin bcd3<=0;bcd2<=9;bcd1<=4;bcd0<=5; end
			946: begin bcd3<=0;bcd2<=9;bcd1<=4;bcd0<=6; end
			947: begin bcd3<=0;bcd2<=9;bcd1<=4;bcd0<=7; end
			948: begin bcd3<=0;bcd2<=9;bcd1<=4;bcd0<=8; end
			949: begin bcd3<=0;bcd2<=9;bcd1<=4;bcd0<=9; end
			950: begin bcd3<=0;bcd2<=9;bcd1<=5;bcd0<=0; end
			951: begin bcd3<=0;bcd2<=9;bcd1<=5;bcd0<=1; end
			952: begin bcd3<=0;bcd2<=9;bcd1<=5;bcd0<=2; end
			953: begin bcd3<=0;bcd2<=9;bcd1<=5;bcd0<=3; end
			954: begin bcd3<=0;bcd2<=9;bcd1<=5;bcd0<=4; end
			955: begin bcd3<=0;bcd2<=9;bcd1<=5;bcd0<=5; end
			956: begin bcd3<=0;bcd2<=9;bcd1<=5;bcd0<=6; end
			957: begin bcd3<=0;bcd2<=9;bcd1<=5;bcd0<=7; end
			958: begin bcd3<=0;bcd2<=9;bcd1<=5;bcd0<=8; end
			959: begin bcd3<=0;bcd2<=9;bcd1<=5;bcd0<=9; end
			960: begin bcd3<=0;bcd2<=9;bcd1<=6;bcd0<=0; end
			961: begin bcd3<=0;bcd2<=9;bcd1<=6;bcd0<=1; end
			962: begin bcd3<=0;bcd2<=9;bcd1<=6;bcd0<=2; end
			963: begin bcd3<=0;bcd2<=9;bcd1<=6;bcd0<=3; end
			964: begin bcd3<=0;bcd2<=9;bcd1<=6;bcd0<=4; end
			965: begin bcd3<=0;bcd2<=9;bcd1<=6;bcd0<=5; end
			966: begin bcd3<=0;bcd2<=9;bcd1<=6;bcd0<=6; end
			967: begin bcd3<=0;bcd2<=9;bcd1<=6;bcd0<=7; end
			968: begin bcd3<=0;bcd2<=9;bcd1<=6;bcd0<=8; end
			969: begin bcd3<=0;bcd2<=9;bcd1<=6;bcd0<=9; end
			970: begin bcd3<=0;bcd2<=9;bcd1<=7;bcd0<=0; end
			971: begin bcd3<=0;bcd2<=9;bcd1<=7;bcd0<=1; end
			972: begin bcd3<=0;bcd2<=9;bcd1<=7;bcd0<=2; end
			973: begin bcd3<=0;bcd2<=9;bcd1<=7;bcd0<=3; end
			974: begin bcd3<=0;bcd2<=9;bcd1<=7;bcd0<=4; end
			975: begin bcd3<=0;bcd2<=9;bcd1<=7;bcd0<=5; end
			976: begin bcd3<=0;bcd2<=9;bcd1<=7;bcd0<=6; end
			977: begin bcd3<=0;bcd2<=9;bcd1<=7;bcd0<=7; end
			978: begin bcd3<=0;bcd2<=9;bcd1<=7;bcd0<=8; end
			979: begin bcd3<=0;bcd2<=9;bcd1<=7;bcd0<=9; end
			980: begin bcd3<=0;bcd2<=9;bcd1<=8;bcd0<=0; end
			981: begin bcd3<=0;bcd2<=9;bcd1<=8;bcd0<=1; end
			982: begin bcd3<=0;bcd2<=9;bcd1<=8;bcd0<=2; end
			983: begin bcd3<=0;bcd2<=9;bcd1<=8;bcd0<=3; end
			984: begin bcd3<=0;bcd2<=9;bcd1<=8;bcd0<=4; end
			985: begin bcd3<=0;bcd2<=9;bcd1<=8;bcd0<=5; end
			986: begin bcd3<=0;bcd2<=9;bcd1<=8;bcd0<=6; end
			987: begin bcd3<=0;bcd2<=9;bcd1<=8;bcd0<=7; end
			988: begin bcd3<=0;bcd2<=9;bcd1<=8;bcd0<=8; end
			989: begin bcd3<=0;bcd2<=9;bcd1<=8;bcd0<=9; end
			990: begin bcd3<=0;bcd2<=9;bcd1<=9;bcd0<=0; end
			991: begin bcd3<=0;bcd2<=9;bcd1<=9;bcd0<=1; end
			992: begin bcd3<=0;bcd2<=9;bcd1<=9;bcd0<=2; end
			993: begin bcd3<=0;bcd2<=9;bcd1<=9;bcd0<=3; end
			994: begin bcd3<=0;bcd2<=9;bcd1<=9;bcd0<=4; end
			995: begin bcd3<=0;bcd2<=9;bcd1<=9;bcd0<=5; end
			996: begin bcd3<=0;bcd2<=9;bcd1<=9;bcd0<=6; end
			997: begin bcd3<=0;bcd2<=9;bcd1<=9;bcd0<=7; end
			998: begin bcd3<=0;bcd2<=9;bcd1<=9;bcd0<=8; end
			999: begin bcd3<=0;bcd2<=9;bcd1<=9;bcd0<=9; end
			1000: begin bcd3<=1;bcd2<=0;bcd1<=0;bcd0<=0; end
			1001: begin bcd3<=1;bcd2<=0;bcd1<=0;bcd0<=1; end
			1002: begin bcd3<=1;bcd2<=0;bcd1<=0;bcd0<=2; end
			1003: begin bcd3<=1;bcd2<=0;bcd1<=0;bcd0<=3; end
			1004: begin bcd3<=1;bcd2<=0;bcd1<=0;bcd0<=4; end
			1005: begin bcd3<=1;bcd2<=0;bcd1<=0;bcd0<=5; end
			1006: begin bcd3<=1;bcd2<=0;bcd1<=0;bcd0<=6; end
			1007: begin bcd3<=1;bcd2<=0;bcd1<=0;bcd0<=7; end
			1008: begin bcd3<=1;bcd2<=0;bcd1<=0;bcd0<=8; end
			1009: begin bcd3<=1;bcd2<=0;bcd1<=0;bcd0<=9; end
			1010: begin bcd3<=1;bcd2<=0;bcd1<=1;bcd0<=0; end
			1011: begin bcd3<=1;bcd2<=0;bcd1<=1;bcd0<=1; end
			1012: begin bcd3<=1;bcd2<=0;bcd1<=1;bcd0<=2; end
			1013: begin bcd3<=1;bcd2<=0;bcd1<=1;bcd0<=3; end
			1014: begin bcd3<=1;bcd2<=0;bcd1<=1;bcd0<=4; end
			1015: begin bcd3<=1;bcd2<=0;bcd1<=1;bcd0<=5; end
			1016: begin bcd3<=1;bcd2<=0;bcd1<=1;bcd0<=6; end
			1017: begin bcd3<=1;bcd2<=0;bcd1<=1;bcd0<=7; end
			1018: begin bcd3<=1;bcd2<=0;bcd1<=1;bcd0<=8; end
			1019: begin bcd3<=1;bcd2<=0;bcd1<=1;bcd0<=9; end
			1020: begin bcd3<=1;bcd2<=0;bcd1<=2;bcd0<=0; end
			1021: begin bcd3<=1;bcd2<=0;bcd1<=2;bcd0<=1; end
			1022: begin bcd3<=1;bcd2<=0;bcd1<=2;bcd0<=2; end
			1023: begin bcd3<=1;bcd2<=0;bcd1<=2;bcd0<=3; end
			1024: begin bcd3<=1;bcd2<=0;bcd1<=2;bcd0<=4; end
			1025: begin bcd3<=1;bcd2<=0;bcd1<=2;bcd0<=5; end
			1026: begin bcd3<=1;bcd2<=0;bcd1<=2;bcd0<=6; end
			1027: begin bcd3<=1;bcd2<=0;bcd1<=2;bcd0<=7; end
			1028: begin bcd3<=1;bcd2<=0;bcd1<=2;bcd0<=8; end
			1029: begin bcd3<=1;bcd2<=0;bcd1<=2;bcd0<=9; end
			1030: begin bcd3<=1;bcd2<=0;bcd1<=3;bcd0<=0; end
			1031: begin bcd3<=1;bcd2<=0;bcd1<=3;bcd0<=1; end
			1032: begin bcd3<=1;bcd2<=0;bcd1<=3;bcd0<=2; end
			1033: begin bcd3<=1;bcd2<=0;bcd1<=3;bcd0<=3; end
			1034: begin bcd3<=1;bcd2<=0;bcd1<=3;bcd0<=4; end
			1035: begin bcd3<=1;bcd2<=0;bcd1<=3;bcd0<=5; end
			1036: begin bcd3<=1;bcd2<=0;bcd1<=3;bcd0<=6; end
			1037: begin bcd3<=1;bcd2<=0;bcd1<=3;bcd0<=7; end
			1038: begin bcd3<=1;bcd2<=0;bcd1<=3;bcd0<=8; end
			1039: begin bcd3<=1;bcd2<=0;bcd1<=3;bcd0<=9; end
			1040: begin bcd3<=1;bcd2<=0;bcd1<=4;bcd0<=0; end
			1041: begin bcd3<=1;bcd2<=0;bcd1<=4;bcd0<=1; end
			1042: begin bcd3<=1;bcd2<=0;bcd1<=4;bcd0<=2; end
			1043: begin bcd3<=1;bcd2<=0;bcd1<=4;bcd0<=3; end
			1044: begin bcd3<=1;bcd2<=0;bcd1<=4;bcd0<=4; end
			1045: begin bcd3<=1;bcd2<=0;bcd1<=4;bcd0<=5; end
			1046: begin bcd3<=1;bcd2<=0;bcd1<=4;bcd0<=6; end
			1047: begin bcd3<=1;bcd2<=0;bcd1<=4;bcd0<=7; end
			1048: begin bcd3<=1;bcd2<=0;bcd1<=4;bcd0<=8; end
			1049: begin bcd3<=1;bcd2<=0;bcd1<=4;bcd0<=9; end
			1050: begin bcd3<=1;bcd2<=0;bcd1<=5;bcd0<=0; end
			1051: begin bcd3<=1;bcd2<=0;bcd1<=5;bcd0<=1; end
			1052: begin bcd3<=1;bcd2<=0;bcd1<=5;bcd0<=2; end
			1053: begin bcd3<=1;bcd2<=0;bcd1<=5;bcd0<=3; end
			1054: begin bcd3<=1;bcd2<=0;bcd1<=5;bcd0<=4; end
			1055: begin bcd3<=1;bcd2<=0;bcd1<=5;bcd0<=5; end
			1056: begin bcd3<=1;bcd2<=0;bcd1<=5;bcd0<=6; end
			1057: begin bcd3<=1;bcd2<=0;bcd1<=5;bcd0<=7; end
			1058: begin bcd3<=1;bcd2<=0;bcd1<=5;bcd0<=8; end
			1059: begin bcd3<=1;bcd2<=0;bcd1<=5;bcd0<=9; end
			1060: begin bcd3<=1;bcd2<=0;bcd1<=6;bcd0<=0; end
			1061: begin bcd3<=1;bcd2<=0;bcd1<=6;bcd0<=1; end
			1062: begin bcd3<=1;bcd2<=0;bcd1<=6;bcd0<=2; end
			1063: begin bcd3<=1;bcd2<=0;bcd1<=6;bcd0<=3; end
			1064: begin bcd3<=1;bcd2<=0;bcd1<=6;bcd0<=4; end
			1065: begin bcd3<=1;bcd2<=0;bcd1<=6;bcd0<=5; end
			1066: begin bcd3<=1;bcd2<=0;bcd1<=6;bcd0<=6; end
			1067: begin bcd3<=1;bcd2<=0;bcd1<=6;bcd0<=7; end
			1068: begin bcd3<=1;bcd2<=0;bcd1<=6;bcd0<=8; end
			1069: begin bcd3<=1;bcd2<=0;bcd1<=6;bcd0<=9; end
			1070: begin bcd3<=1;bcd2<=0;bcd1<=7;bcd0<=0; end
			1071: begin bcd3<=1;bcd2<=0;bcd1<=7;bcd0<=1; end
			1072: begin bcd3<=1;bcd2<=0;bcd1<=7;bcd0<=2; end
			1073: begin bcd3<=1;bcd2<=0;bcd1<=7;bcd0<=3; end
			1074: begin bcd3<=1;bcd2<=0;bcd1<=7;bcd0<=4; end
			1075: begin bcd3<=1;bcd2<=0;bcd1<=7;bcd0<=5; end
			1076: begin bcd3<=1;bcd2<=0;bcd1<=7;bcd0<=6; end
			1077: begin bcd3<=1;bcd2<=0;bcd1<=7;bcd0<=7; end
			1078: begin bcd3<=1;bcd2<=0;bcd1<=7;bcd0<=8; end
			1079: begin bcd3<=1;bcd2<=0;bcd1<=7;bcd0<=9; end
			1080: begin bcd3<=1;bcd2<=0;bcd1<=8;bcd0<=0; end
			1081: begin bcd3<=1;bcd2<=0;bcd1<=8;bcd0<=1; end
			1082: begin bcd3<=1;bcd2<=0;bcd1<=8;bcd0<=2; end
			1083: begin bcd3<=1;bcd2<=0;bcd1<=8;bcd0<=3; end
			1084: begin bcd3<=1;bcd2<=0;bcd1<=8;bcd0<=4; end
			1085: begin bcd3<=1;bcd2<=0;bcd1<=8;bcd0<=5; end
			1086: begin bcd3<=1;bcd2<=0;bcd1<=8;bcd0<=6; end
			1087: begin bcd3<=1;bcd2<=0;bcd1<=8;bcd0<=7; end
			1088: begin bcd3<=1;bcd2<=0;bcd1<=8;bcd0<=8; end
			1089: begin bcd3<=1;bcd2<=0;bcd1<=8;bcd0<=9; end
			1090: begin bcd3<=1;bcd2<=0;bcd1<=9;bcd0<=0; end
			1091: begin bcd3<=1;bcd2<=0;bcd1<=9;bcd0<=1; end
			1092: begin bcd3<=1;bcd2<=0;bcd1<=9;bcd0<=2; end
			1093: begin bcd3<=1;bcd2<=0;bcd1<=9;bcd0<=3; end
			1094: begin bcd3<=1;bcd2<=0;bcd1<=9;bcd0<=4; end
			1095: begin bcd3<=1;bcd2<=0;bcd1<=9;bcd0<=5; end
			1096: begin bcd3<=1;bcd2<=0;bcd1<=9;bcd0<=6; end
			1097: begin bcd3<=1;bcd2<=0;bcd1<=9;bcd0<=7; end
			1098: begin bcd3<=1;bcd2<=0;bcd1<=9;bcd0<=8; end
			1099: begin bcd3<=1;bcd2<=0;bcd1<=9;bcd0<=9; end
			1100: begin bcd3<=1;bcd2<=1;bcd1<=0;bcd0<=0; end
			1101: begin bcd3<=1;bcd2<=1;bcd1<=0;bcd0<=1; end
			1102: begin bcd3<=1;bcd2<=1;bcd1<=0;bcd0<=2; end
			1103: begin bcd3<=1;bcd2<=1;bcd1<=0;bcd0<=3; end
			1104: begin bcd3<=1;bcd2<=1;bcd1<=0;bcd0<=4; end
			1105: begin bcd3<=1;bcd2<=1;bcd1<=0;bcd0<=5; end
			1106: begin bcd3<=1;bcd2<=1;bcd1<=0;bcd0<=6; end
			1107: begin bcd3<=1;bcd2<=1;bcd1<=0;bcd0<=7; end
			1108: begin bcd3<=1;bcd2<=1;bcd1<=0;bcd0<=8; end
			1109: begin bcd3<=1;bcd2<=1;bcd1<=0;bcd0<=9; end
			1110: begin bcd3<=1;bcd2<=1;bcd1<=1;bcd0<=0; end
			1111: begin bcd3<=1;bcd2<=1;bcd1<=1;bcd0<=1; end
			1112: begin bcd3<=1;bcd2<=1;bcd1<=1;bcd0<=2; end
			1113: begin bcd3<=1;bcd2<=1;bcd1<=1;bcd0<=3; end
			1114: begin bcd3<=1;bcd2<=1;bcd1<=1;bcd0<=4; end
			1115: begin bcd3<=1;bcd2<=1;bcd1<=1;bcd0<=5; end
			1116: begin bcd3<=1;bcd2<=1;bcd1<=1;bcd0<=6; end
			1117: begin bcd3<=1;bcd2<=1;bcd1<=1;bcd0<=7; end
			1118: begin bcd3<=1;bcd2<=1;bcd1<=1;bcd0<=8; end
			1119: begin bcd3<=1;bcd2<=1;bcd1<=1;bcd0<=9; end
			1120: begin bcd3<=1;bcd2<=1;bcd1<=2;bcd0<=0; end
			1121: begin bcd3<=1;bcd2<=1;bcd1<=2;bcd0<=1; end
			1122: begin bcd3<=1;bcd2<=1;bcd1<=2;bcd0<=2; end
			1123: begin bcd3<=1;bcd2<=1;bcd1<=2;bcd0<=3; end
			1124: begin bcd3<=1;bcd2<=1;bcd1<=2;bcd0<=4; end
			1125: begin bcd3<=1;bcd2<=1;bcd1<=2;bcd0<=5; end
			1126: begin bcd3<=1;bcd2<=1;bcd1<=2;bcd0<=6; end
			1127: begin bcd3<=1;bcd2<=1;bcd1<=2;bcd0<=7; end
			1128: begin bcd3<=1;bcd2<=1;bcd1<=2;bcd0<=8; end
			1129: begin bcd3<=1;bcd2<=1;bcd1<=2;bcd0<=9; end
			1130: begin bcd3<=1;bcd2<=1;bcd1<=3;bcd0<=0; end
			1131: begin bcd3<=1;bcd2<=1;bcd1<=3;bcd0<=1; end
			1132: begin bcd3<=1;bcd2<=1;bcd1<=3;bcd0<=2; end
			1133: begin bcd3<=1;bcd2<=1;bcd1<=3;bcd0<=3; end
			1134: begin bcd3<=1;bcd2<=1;bcd1<=3;bcd0<=4; end
			1135: begin bcd3<=1;bcd2<=1;bcd1<=3;bcd0<=5; end
			1136: begin bcd3<=1;bcd2<=1;bcd1<=3;bcd0<=6; end
			1137: begin bcd3<=1;bcd2<=1;bcd1<=3;bcd0<=7; end
			1138: begin bcd3<=1;bcd2<=1;bcd1<=3;bcd0<=8; end
			1139: begin bcd3<=1;bcd2<=1;bcd1<=3;bcd0<=9; end
			1140: begin bcd3<=1;bcd2<=1;bcd1<=4;bcd0<=0; end
			1141: begin bcd3<=1;bcd2<=1;bcd1<=4;bcd0<=1; end
			1142: begin bcd3<=1;bcd2<=1;bcd1<=4;bcd0<=2; end
			1143: begin bcd3<=1;bcd2<=1;bcd1<=4;bcd0<=3; end
			1144: begin bcd3<=1;bcd2<=1;bcd1<=4;bcd0<=4; end
			1145: begin bcd3<=1;bcd2<=1;bcd1<=4;bcd0<=5; end
			1146: begin bcd3<=1;bcd2<=1;bcd1<=4;bcd0<=6; end
			1147: begin bcd3<=1;bcd2<=1;bcd1<=4;bcd0<=7; end
			1148: begin bcd3<=1;bcd2<=1;bcd1<=4;bcd0<=8; end
			1149: begin bcd3<=1;bcd2<=1;bcd1<=4;bcd0<=9; end
			1150: begin bcd3<=1;bcd2<=1;bcd1<=5;bcd0<=0; end
			1151: begin bcd3<=1;bcd2<=1;bcd1<=5;bcd0<=1; end
			1152: begin bcd3<=1;bcd2<=1;bcd1<=5;bcd0<=2; end
			1153: begin bcd3<=1;bcd2<=1;bcd1<=5;bcd0<=3; end
			1154: begin bcd3<=1;bcd2<=1;bcd1<=5;bcd0<=4; end
			1155: begin bcd3<=1;bcd2<=1;bcd1<=5;bcd0<=5; end
			1156: begin bcd3<=1;bcd2<=1;bcd1<=5;bcd0<=6; end
			1157: begin bcd3<=1;bcd2<=1;bcd1<=5;bcd0<=7; end
			1158: begin bcd3<=1;bcd2<=1;bcd1<=5;bcd0<=8; end
			1159: begin bcd3<=1;bcd2<=1;bcd1<=5;bcd0<=9; end
			1160: begin bcd3<=1;bcd2<=1;bcd1<=6;bcd0<=0; end
			1161: begin bcd3<=1;bcd2<=1;bcd1<=6;bcd0<=1; end
			1162: begin bcd3<=1;bcd2<=1;bcd1<=6;bcd0<=2; end
			1163: begin bcd3<=1;bcd2<=1;bcd1<=6;bcd0<=3; end
			1164: begin bcd3<=1;bcd2<=1;bcd1<=6;bcd0<=4; end
			1165: begin bcd3<=1;bcd2<=1;bcd1<=6;bcd0<=5; end
			1166: begin bcd3<=1;bcd2<=1;bcd1<=6;bcd0<=6; end
			1167: begin bcd3<=1;bcd2<=1;bcd1<=6;bcd0<=7; end
			1168: begin bcd3<=1;bcd2<=1;bcd1<=6;bcd0<=8; end
			1169: begin bcd3<=1;bcd2<=1;bcd1<=6;bcd0<=9; end
			1170: begin bcd3<=1;bcd2<=1;bcd1<=7;bcd0<=0; end
			1171: begin bcd3<=1;bcd2<=1;bcd1<=7;bcd0<=1; end
			1172: begin bcd3<=1;bcd2<=1;bcd1<=7;bcd0<=2; end
			1173: begin bcd3<=1;bcd2<=1;bcd1<=7;bcd0<=3; end
			1174: begin bcd3<=1;bcd2<=1;bcd1<=7;bcd0<=4; end
			1175: begin bcd3<=1;bcd2<=1;bcd1<=7;bcd0<=5; end
			1176: begin bcd3<=1;bcd2<=1;bcd1<=7;bcd0<=6; end
			1177: begin bcd3<=1;bcd2<=1;bcd1<=7;bcd0<=7; end
			1178: begin bcd3<=1;bcd2<=1;bcd1<=7;bcd0<=8; end
			1179: begin bcd3<=1;bcd2<=1;bcd1<=7;bcd0<=9; end
			1180: begin bcd3<=1;bcd2<=1;bcd1<=8;bcd0<=0; end
			1181: begin bcd3<=1;bcd2<=1;bcd1<=8;bcd0<=1; end
			1182: begin bcd3<=1;bcd2<=1;bcd1<=8;bcd0<=2; end
			1183: begin bcd3<=1;bcd2<=1;bcd1<=8;bcd0<=3; end
			1184: begin bcd3<=1;bcd2<=1;bcd1<=8;bcd0<=4; end
			1185: begin bcd3<=1;bcd2<=1;bcd1<=8;bcd0<=5; end
			1186: begin bcd3<=1;bcd2<=1;bcd1<=8;bcd0<=6; end
			1187: begin bcd3<=1;bcd2<=1;bcd1<=8;bcd0<=7; end
			1188: begin bcd3<=1;bcd2<=1;bcd1<=8;bcd0<=8; end
			1189: begin bcd3<=1;bcd2<=1;bcd1<=8;bcd0<=9; end
			1190: begin bcd3<=1;bcd2<=1;bcd1<=9;bcd0<=0; end
			1191: begin bcd3<=1;bcd2<=1;bcd1<=9;bcd0<=1; end
			1192: begin bcd3<=1;bcd2<=1;bcd1<=9;bcd0<=2; end
			1193: begin bcd3<=1;bcd2<=1;bcd1<=9;bcd0<=3; end
			1194: begin bcd3<=1;bcd2<=1;bcd1<=9;bcd0<=4; end
			1195: begin bcd3<=1;bcd2<=1;bcd1<=9;bcd0<=5; end
			1196: begin bcd3<=1;bcd2<=1;bcd1<=9;bcd0<=6; end
			1197: begin bcd3<=1;bcd2<=1;bcd1<=9;bcd0<=7; end
			1198: begin bcd3<=1;bcd2<=1;bcd1<=9;bcd0<=8; end
			1199: begin bcd3<=1;bcd2<=1;bcd1<=9;bcd0<=9; end
			1200: begin bcd3<=1;bcd2<=2;bcd1<=0;bcd0<=0; end
			1201: begin bcd3<=1;bcd2<=2;bcd1<=0;bcd0<=1; end
			1202: begin bcd3<=1;bcd2<=2;bcd1<=0;bcd0<=2; end
			1203: begin bcd3<=1;bcd2<=2;bcd1<=0;bcd0<=3; end
			1204: begin bcd3<=1;bcd2<=2;bcd1<=0;bcd0<=4; end
			1205: begin bcd3<=1;bcd2<=2;bcd1<=0;bcd0<=5; end
			1206: begin bcd3<=1;bcd2<=2;bcd1<=0;bcd0<=6; end
			1207: begin bcd3<=1;bcd2<=2;bcd1<=0;bcd0<=7; end
			1208: begin bcd3<=1;bcd2<=2;bcd1<=0;bcd0<=8; end
			1209: begin bcd3<=1;bcd2<=2;bcd1<=0;bcd0<=9; end
			1210: begin bcd3<=1;bcd2<=2;bcd1<=1;bcd0<=0; end
			1211: begin bcd3<=1;bcd2<=2;bcd1<=1;bcd0<=1; end
			1212: begin bcd3<=1;bcd2<=2;bcd1<=1;bcd0<=2; end
			1213: begin bcd3<=1;bcd2<=2;bcd1<=1;bcd0<=3; end
			1214: begin bcd3<=1;bcd2<=2;bcd1<=1;bcd0<=4; end
			1215: begin bcd3<=1;bcd2<=2;bcd1<=1;bcd0<=5; end
			1216: begin bcd3<=1;bcd2<=2;bcd1<=1;bcd0<=6; end
			1217: begin bcd3<=1;bcd2<=2;bcd1<=1;bcd0<=7; end
			1218: begin bcd3<=1;bcd2<=2;bcd1<=1;bcd0<=8; end
			1219: begin bcd3<=1;bcd2<=2;bcd1<=1;bcd0<=9; end
			1220: begin bcd3<=1;bcd2<=2;bcd1<=2;bcd0<=0; end
			1221: begin bcd3<=1;bcd2<=2;bcd1<=2;bcd0<=1; end
			1222: begin bcd3<=1;bcd2<=2;bcd1<=2;bcd0<=2; end
			1223: begin bcd3<=1;bcd2<=2;bcd1<=2;bcd0<=3; end
			1224: begin bcd3<=1;bcd2<=2;bcd1<=2;bcd0<=4; end
			1225: begin bcd3<=1;bcd2<=2;bcd1<=2;bcd0<=5; end
			1226: begin bcd3<=1;bcd2<=2;bcd1<=2;bcd0<=6; end
			1227: begin bcd3<=1;bcd2<=2;bcd1<=2;bcd0<=7; end
			1228: begin bcd3<=1;bcd2<=2;bcd1<=2;bcd0<=8; end
			1229: begin bcd3<=1;bcd2<=2;bcd1<=2;bcd0<=9; end
			1230: begin bcd3<=1;bcd2<=2;bcd1<=3;bcd0<=0; end
			1231: begin bcd3<=1;bcd2<=2;bcd1<=3;bcd0<=1; end
			1232: begin bcd3<=1;bcd2<=2;bcd1<=3;bcd0<=2; end
			1233: begin bcd3<=1;bcd2<=2;bcd1<=3;bcd0<=3; end
			1234: begin bcd3<=1;bcd2<=2;bcd1<=3;bcd0<=4; end
			1235: begin bcd3<=1;bcd2<=2;bcd1<=3;bcd0<=5; end
			1236: begin bcd3<=1;bcd2<=2;bcd1<=3;bcd0<=6; end
			1237: begin bcd3<=1;bcd2<=2;bcd1<=3;bcd0<=7; end
			1238: begin bcd3<=1;bcd2<=2;bcd1<=3;bcd0<=8; end
			1239: begin bcd3<=1;bcd2<=2;bcd1<=3;bcd0<=9; end
			1240: begin bcd3<=1;bcd2<=2;bcd1<=4;bcd0<=0; end
			1241: begin bcd3<=1;bcd2<=2;bcd1<=4;bcd0<=1; end
			1242: begin bcd3<=1;bcd2<=2;bcd1<=4;bcd0<=2; end
			1243: begin bcd3<=1;bcd2<=2;bcd1<=4;bcd0<=3; end
			1244: begin bcd3<=1;bcd2<=2;bcd1<=4;bcd0<=4; end
			1245: begin bcd3<=1;bcd2<=2;bcd1<=4;bcd0<=5; end
			1246: begin bcd3<=1;bcd2<=2;bcd1<=4;bcd0<=6; end
			1247: begin bcd3<=1;bcd2<=2;bcd1<=4;bcd0<=7; end
			1248: begin bcd3<=1;bcd2<=2;bcd1<=4;bcd0<=8; end
			1249: begin bcd3<=1;bcd2<=2;bcd1<=4;bcd0<=9; end
			1250: begin bcd3<=1;bcd2<=2;bcd1<=5;bcd0<=0; end
			1251: begin bcd3<=1;bcd2<=2;bcd1<=5;bcd0<=1; end
			1252: begin bcd3<=1;bcd2<=2;bcd1<=5;bcd0<=2; end
			1253: begin bcd3<=1;bcd2<=2;bcd1<=5;bcd0<=3; end
			1254: begin bcd3<=1;bcd2<=2;bcd1<=5;bcd0<=4; end
			1255: begin bcd3<=1;bcd2<=2;bcd1<=5;bcd0<=5; end
			1256: begin bcd3<=1;bcd2<=2;bcd1<=5;bcd0<=6; end
			1257: begin bcd3<=1;bcd2<=2;bcd1<=5;bcd0<=7; end
			1258: begin bcd3<=1;bcd2<=2;bcd1<=5;bcd0<=8; end
			1259: begin bcd3<=1;bcd2<=2;bcd1<=5;bcd0<=9; end
			1260: begin bcd3<=1;bcd2<=2;bcd1<=6;bcd0<=0; end
			1261: begin bcd3<=1;bcd2<=2;bcd1<=6;bcd0<=1; end
			1262: begin bcd3<=1;bcd2<=2;bcd1<=6;bcd0<=2; end
			1263: begin bcd3<=1;bcd2<=2;bcd1<=6;bcd0<=3; end
			1264: begin bcd3<=1;bcd2<=2;bcd1<=6;bcd0<=4; end
			1265: begin bcd3<=1;bcd2<=2;bcd1<=6;bcd0<=5; end
			1266: begin bcd3<=1;bcd2<=2;bcd1<=6;bcd0<=6; end
			1267: begin bcd3<=1;bcd2<=2;bcd1<=6;bcd0<=7; end
			1268: begin bcd3<=1;bcd2<=2;bcd1<=6;bcd0<=8; end
			1269: begin bcd3<=1;bcd2<=2;bcd1<=6;bcd0<=9; end
			1270: begin bcd3<=1;bcd2<=2;bcd1<=7;bcd0<=0; end
			1271: begin bcd3<=1;bcd2<=2;bcd1<=7;bcd0<=1; end
			1272: begin bcd3<=1;bcd2<=2;bcd1<=7;bcd0<=2; end
			1273: begin bcd3<=1;bcd2<=2;bcd1<=7;bcd0<=3; end
			1274: begin bcd3<=1;bcd2<=2;bcd1<=7;bcd0<=4; end
			1275: begin bcd3<=1;bcd2<=2;bcd1<=7;bcd0<=5; end
			1276: begin bcd3<=1;bcd2<=2;bcd1<=7;bcd0<=6; end
			1277: begin bcd3<=1;bcd2<=2;bcd1<=7;bcd0<=7; end
			1278: begin bcd3<=1;bcd2<=2;bcd1<=7;bcd0<=8; end
			1279: begin bcd3<=1;bcd2<=2;bcd1<=7;bcd0<=9; end
			1280: begin bcd3<=1;bcd2<=2;bcd1<=8;bcd0<=0; end
			1281: begin bcd3<=1;bcd2<=2;bcd1<=8;bcd0<=1; end
			1282: begin bcd3<=1;bcd2<=2;bcd1<=8;bcd0<=2; end
			1283: begin bcd3<=1;bcd2<=2;bcd1<=8;bcd0<=3; end
			1284: begin bcd3<=1;bcd2<=2;bcd1<=8;bcd0<=4; end
			1285: begin bcd3<=1;bcd2<=2;bcd1<=8;bcd0<=5; end
			1286: begin bcd3<=1;bcd2<=2;bcd1<=8;bcd0<=6; end
			1287: begin bcd3<=1;bcd2<=2;bcd1<=8;bcd0<=7; end
			1288: begin bcd3<=1;bcd2<=2;bcd1<=8;bcd0<=8; end
			1289: begin bcd3<=1;bcd2<=2;bcd1<=8;bcd0<=9; end
			1290: begin bcd3<=1;bcd2<=2;bcd1<=9;bcd0<=0; end
			1291: begin bcd3<=1;bcd2<=2;bcd1<=9;bcd0<=1; end
			1292: begin bcd3<=1;bcd2<=2;bcd1<=9;bcd0<=2; end
			1293: begin bcd3<=1;bcd2<=2;bcd1<=9;bcd0<=3; end
			1294: begin bcd3<=1;bcd2<=2;bcd1<=9;bcd0<=4; end
			1295: begin bcd3<=1;bcd2<=2;bcd1<=9;bcd0<=5; end
			1296: begin bcd3<=1;bcd2<=2;bcd1<=9;bcd0<=6; end
			1297: begin bcd3<=1;bcd2<=2;bcd1<=9;bcd0<=7; end
			1298: begin bcd3<=1;bcd2<=2;bcd1<=9;bcd0<=8; end
			1299: begin bcd3<=1;bcd2<=2;bcd1<=9;bcd0<=9; end
			1300: begin bcd3<=1;bcd2<=3;bcd1<=0;bcd0<=0; end
			1301: begin bcd3<=1;bcd2<=3;bcd1<=0;bcd0<=1; end
			1302: begin bcd3<=1;bcd2<=3;bcd1<=0;bcd0<=2; end
			1303: begin bcd3<=1;bcd2<=3;bcd1<=0;bcd0<=3; end
			1304: begin bcd3<=1;bcd2<=3;bcd1<=0;bcd0<=4; end
			1305: begin bcd3<=1;bcd2<=3;bcd1<=0;bcd0<=5; end
			1306: begin bcd3<=1;bcd2<=3;bcd1<=0;bcd0<=6; end
			1307: begin bcd3<=1;bcd2<=3;bcd1<=0;bcd0<=7; end
			1308: begin bcd3<=1;bcd2<=3;bcd1<=0;bcd0<=8; end
			1309: begin bcd3<=1;bcd2<=3;bcd1<=0;bcd0<=9; end
			1310: begin bcd3<=1;bcd2<=3;bcd1<=1;bcd0<=0; end
			1311: begin bcd3<=1;bcd2<=3;bcd1<=1;bcd0<=1; end
			1312: begin bcd3<=1;bcd2<=3;bcd1<=1;bcd0<=2; end
			1313: begin bcd3<=1;bcd2<=3;bcd1<=1;bcd0<=3; end
			1314: begin bcd3<=1;bcd2<=3;bcd1<=1;bcd0<=4; end
			1315: begin bcd3<=1;bcd2<=3;bcd1<=1;bcd0<=5; end
			1316: begin bcd3<=1;bcd2<=3;bcd1<=1;bcd0<=6; end
			1317: begin bcd3<=1;bcd2<=3;bcd1<=1;bcd0<=7; end
			1318: begin bcd3<=1;bcd2<=3;bcd1<=1;bcd0<=8; end
			1319: begin bcd3<=1;bcd2<=3;bcd1<=1;bcd0<=9; end
			1320: begin bcd3<=1;bcd2<=3;bcd1<=2;bcd0<=0; end
			1321: begin bcd3<=1;bcd2<=3;bcd1<=2;bcd0<=1; end
			1322: begin bcd3<=1;bcd2<=3;bcd1<=2;bcd0<=2; end
			1323: begin bcd3<=1;bcd2<=3;bcd1<=2;bcd0<=3; end
			1324: begin bcd3<=1;bcd2<=3;bcd1<=2;bcd0<=4; end
			1325: begin bcd3<=1;bcd2<=3;bcd1<=2;bcd0<=5; end
			1326: begin bcd3<=1;bcd2<=3;bcd1<=2;bcd0<=6; end
			1327: begin bcd3<=1;bcd2<=3;bcd1<=2;bcd0<=7; end
			1328: begin bcd3<=1;bcd2<=3;bcd1<=2;bcd0<=8; end
			1329: begin bcd3<=1;bcd2<=3;bcd1<=2;bcd0<=9; end
			1330: begin bcd3<=1;bcd2<=3;bcd1<=3;bcd0<=0; end
			1331: begin bcd3<=1;bcd2<=3;bcd1<=3;bcd0<=1; end
			1332: begin bcd3<=1;bcd2<=3;bcd1<=3;bcd0<=2; end
			1333: begin bcd3<=1;bcd2<=3;bcd1<=3;bcd0<=3; end
			1334: begin bcd3<=1;bcd2<=3;bcd1<=3;bcd0<=4; end
			1335: begin bcd3<=1;bcd2<=3;bcd1<=3;bcd0<=5; end
			1336: begin bcd3<=1;bcd2<=3;bcd1<=3;bcd0<=6; end
			1337: begin bcd3<=1;bcd2<=3;bcd1<=3;bcd0<=7; end
			1338: begin bcd3<=1;bcd2<=3;bcd1<=3;bcd0<=8; end
			1339: begin bcd3<=1;bcd2<=3;bcd1<=3;bcd0<=9; end
			1340: begin bcd3<=1;bcd2<=3;bcd1<=4;bcd0<=0; end
			1341: begin bcd3<=1;bcd2<=3;bcd1<=4;bcd0<=1; end
			1342: begin bcd3<=1;bcd2<=3;bcd1<=4;bcd0<=2; end
			1343: begin bcd3<=1;bcd2<=3;bcd1<=4;bcd0<=3; end
			1344: begin bcd3<=1;bcd2<=3;bcd1<=4;bcd0<=4; end
			1345: begin bcd3<=1;bcd2<=3;bcd1<=4;bcd0<=5; end
			1346: begin bcd3<=1;bcd2<=3;bcd1<=4;bcd0<=6; end
			1347: begin bcd3<=1;bcd2<=3;bcd1<=4;bcd0<=7; end
			1348: begin bcd3<=1;bcd2<=3;bcd1<=4;bcd0<=8; end
			1349: begin bcd3<=1;bcd2<=3;bcd1<=4;bcd0<=9; end
			1350: begin bcd3<=1;bcd2<=3;bcd1<=5;bcd0<=0; end
			1351: begin bcd3<=1;bcd2<=3;bcd1<=5;bcd0<=1; end
			1352: begin bcd3<=1;bcd2<=3;bcd1<=5;bcd0<=2; end
			1353: begin bcd3<=1;bcd2<=3;bcd1<=5;bcd0<=3; end
			1354: begin bcd3<=1;bcd2<=3;bcd1<=5;bcd0<=4; end
			1355: begin bcd3<=1;bcd2<=3;bcd1<=5;bcd0<=5; end
			1356: begin bcd3<=1;bcd2<=3;bcd1<=5;bcd0<=6; end
			1357: begin bcd3<=1;bcd2<=3;bcd1<=5;bcd0<=7; end
			1358: begin bcd3<=1;bcd2<=3;bcd1<=5;bcd0<=8; end
			1359: begin bcd3<=1;bcd2<=3;bcd1<=5;bcd0<=9; end
			1360: begin bcd3<=1;bcd2<=3;bcd1<=6;bcd0<=0; end
			1361: begin bcd3<=1;bcd2<=3;bcd1<=6;bcd0<=1; end
			1362: begin bcd3<=1;bcd2<=3;bcd1<=6;bcd0<=2; end
			1363: begin bcd3<=1;bcd2<=3;bcd1<=6;bcd0<=3; end
			1364: begin bcd3<=1;bcd2<=3;bcd1<=6;bcd0<=4; end
			1365: begin bcd3<=1;bcd2<=3;bcd1<=6;bcd0<=5; end
			1366: begin bcd3<=1;bcd2<=3;bcd1<=6;bcd0<=6; end
			1367: begin bcd3<=1;bcd2<=3;bcd1<=6;bcd0<=7; end
			1368: begin bcd3<=1;bcd2<=3;bcd1<=6;bcd0<=8; end
			1369: begin bcd3<=1;bcd2<=3;bcd1<=6;bcd0<=9; end
			1370: begin bcd3<=1;bcd2<=3;bcd1<=7;bcd0<=0; end
			1371: begin bcd3<=1;bcd2<=3;bcd1<=7;bcd0<=1; end
			1372: begin bcd3<=1;bcd2<=3;bcd1<=7;bcd0<=2; end
			1373: begin bcd3<=1;bcd2<=3;bcd1<=7;bcd0<=3; end
			1374: begin bcd3<=1;bcd2<=3;bcd1<=7;bcd0<=4; end
			1375: begin bcd3<=1;bcd2<=3;bcd1<=7;bcd0<=5; end
			1376: begin bcd3<=1;bcd2<=3;bcd1<=7;bcd0<=6; end
			1377: begin bcd3<=1;bcd2<=3;bcd1<=7;bcd0<=7; end
			1378: begin bcd3<=1;bcd2<=3;bcd1<=7;bcd0<=8; end
			1379: begin bcd3<=1;bcd2<=3;bcd1<=7;bcd0<=9; end
			1380: begin bcd3<=1;bcd2<=3;bcd1<=8;bcd0<=0; end
			1381: begin bcd3<=1;bcd2<=3;bcd1<=8;bcd0<=1; end
			1382: begin bcd3<=1;bcd2<=3;bcd1<=8;bcd0<=2; end
			1383: begin bcd3<=1;bcd2<=3;bcd1<=8;bcd0<=3; end
			1384: begin bcd3<=1;bcd2<=3;bcd1<=8;bcd0<=4; end
			1385: begin bcd3<=1;bcd2<=3;bcd1<=8;bcd0<=5; end
			1386: begin bcd3<=1;bcd2<=3;bcd1<=8;bcd0<=6; end
			1387: begin bcd3<=1;bcd2<=3;bcd1<=8;bcd0<=7; end
			1388: begin bcd3<=1;bcd2<=3;bcd1<=8;bcd0<=8; end
			1389: begin bcd3<=1;bcd2<=3;bcd1<=8;bcd0<=9; end
			1390: begin bcd3<=1;bcd2<=3;bcd1<=9;bcd0<=0; end
			1391: begin bcd3<=1;bcd2<=3;bcd1<=9;bcd0<=1; end
			1392: begin bcd3<=1;bcd2<=3;bcd1<=9;bcd0<=2; end
			1393: begin bcd3<=1;bcd2<=3;bcd1<=9;bcd0<=3; end
			1394: begin bcd3<=1;bcd2<=3;bcd1<=9;bcd0<=4; end
			1395: begin bcd3<=1;bcd2<=3;bcd1<=9;bcd0<=5; end
			1396: begin bcd3<=1;bcd2<=3;bcd1<=9;bcd0<=6; end
			1397: begin bcd3<=1;bcd2<=3;bcd1<=9;bcd0<=7; end
			1398: begin bcd3<=1;bcd2<=3;bcd1<=9;bcd0<=8; end
			1399: begin bcd3<=1;bcd2<=3;bcd1<=9;bcd0<=9; end
			1400: begin bcd3<=1;bcd2<=4;bcd1<=0;bcd0<=0; end
			1401: begin bcd3<=1;bcd2<=4;bcd1<=0;bcd0<=1; end
			1402: begin bcd3<=1;bcd2<=4;bcd1<=0;bcd0<=2; end
			1403: begin bcd3<=1;bcd2<=4;bcd1<=0;bcd0<=3; end
			1404: begin bcd3<=1;bcd2<=4;bcd1<=0;bcd0<=4; end
			1405: begin bcd3<=1;bcd2<=4;bcd1<=0;bcd0<=5; end
			1406: begin bcd3<=1;bcd2<=4;bcd1<=0;bcd0<=6; end
			1407: begin bcd3<=1;bcd2<=4;bcd1<=0;bcd0<=7; end
			1408: begin bcd3<=1;bcd2<=4;bcd1<=0;bcd0<=8; end
			1409: begin bcd3<=1;bcd2<=4;bcd1<=0;bcd0<=9; end
			1410: begin bcd3<=1;bcd2<=4;bcd1<=1;bcd0<=0; end
			1411: begin bcd3<=1;bcd2<=4;bcd1<=1;bcd0<=1; end
			1412: begin bcd3<=1;bcd2<=4;bcd1<=1;bcd0<=2; end
			1413: begin bcd3<=1;bcd2<=4;bcd1<=1;bcd0<=3; end
			1414: begin bcd3<=1;bcd2<=4;bcd1<=1;bcd0<=4; end
			1415: begin bcd3<=1;bcd2<=4;bcd1<=1;bcd0<=5; end
			1416: begin bcd3<=1;bcd2<=4;bcd1<=1;bcd0<=6; end
			1417: begin bcd3<=1;bcd2<=4;bcd1<=1;bcd0<=7; end
			1418: begin bcd3<=1;bcd2<=4;bcd1<=1;bcd0<=8; end
			1419: begin bcd3<=1;bcd2<=4;bcd1<=1;bcd0<=9; end
			1420: begin bcd3<=1;bcd2<=4;bcd1<=2;bcd0<=0; end
			1421: begin bcd3<=1;bcd2<=4;bcd1<=2;bcd0<=1; end
			1422: begin bcd3<=1;bcd2<=4;bcd1<=2;bcd0<=2; end
			1423: begin bcd3<=1;bcd2<=4;bcd1<=2;bcd0<=3; end
			1424: begin bcd3<=1;bcd2<=4;bcd1<=2;bcd0<=4; end
			1425: begin bcd3<=1;bcd2<=4;bcd1<=2;bcd0<=5; end
			1426: begin bcd3<=1;bcd2<=4;bcd1<=2;bcd0<=6; end
			1427: begin bcd3<=1;bcd2<=4;bcd1<=2;bcd0<=7; end
			1428: begin bcd3<=1;bcd2<=4;bcd1<=2;bcd0<=8; end
			1429: begin bcd3<=1;bcd2<=4;bcd1<=2;bcd0<=9; end
			1430: begin bcd3<=1;bcd2<=4;bcd1<=3;bcd0<=0; end
			1431: begin bcd3<=1;bcd2<=4;bcd1<=3;bcd0<=1; end
			1432: begin bcd3<=1;bcd2<=4;bcd1<=3;bcd0<=2; end
			1433: begin bcd3<=1;bcd2<=4;bcd1<=3;bcd0<=3; end
			1434: begin bcd3<=1;bcd2<=4;bcd1<=3;bcd0<=4; end
			1435: begin bcd3<=1;bcd2<=4;bcd1<=3;bcd0<=5; end
			1436: begin bcd3<=1;bcd2<=4;bcd1<=3;bcd0<=6; end
			1437: begin bcd3<=1;bcd2<=4;bcd1<=3;bcd0<=7; end
			1438: begin bcd3<=1;bcd2<=4;bcd1<=3;bcd0<=8; end
			1439: begin bcd3<=1;bcd2<=4;bcd1<=3;bcd0<=9; end
			1440: begin bcd3<=1;bcd2<=4;bcd1<=4;bcd0<=0; end
			1441: begin bcd3<=1;bcd2<=4;bcd1<=4;bcd0<=1; end
			1442: begin bcd3<=1;bcd2<=4;bcd1<=4;bcd0<=2; end
			1443: begin bcd3<=1;bcd2<=4;bcd1<=4;bcd0<=3; end
			1444: begin bcd3<=1;bcd2<=4;bcd1<=4;bcd0<=4; end
			1445: begin bcd3<=1;bcd2<=4;bcd1<=4;bcd0<=5; end
			1446: begin bcd3<=1;bcd2<=4;bcd1<=4;bcd0<=6; end
			1447: begin bcd3<=1;bcd2<=4;bcd1<=4;bcd0<=7; end
			1448: begin bcd3<=1;bcd2<=4;bcd1<=4;bcd0<=8; end
			1449: begin bcd3<=1;bcd2<=4;bcd1<=4;bcd0<=9; end
			1450: begin bcd3<=1;bcd2<=4;bcd1<=5;bcd0<=0; end
			1451: begin bcd3<=1;bcd2<=4;bcd1<=5;bcd0<=1; end
			1452: begin bcd3<=1;bcd2<=4;bcd1<=5;bcd0<=2; end
			1453: begin bcd3<=1;bcd2<=4;bcd1<=5;bcd0<=3; end
			1454: begin bcd3<=1;bcd2<=4;bcd1<=5;bcd0<=4; end
			1455: begin bcd3<=1;bcd2<=4;bcd1<=5;bcd0<=5; end
			1456: begin bcd3<=1;bcd2<=4;bcd1<=5;bcd0<=6; end
			1457: begin bcd3<=1;bcd2<=4;bcd1<=5;bcd0<=7; end
			1458: begin bcd3<=1;bcd2<=4;bcd1<=5;bcd0<=8; end
			1459: begin bcd3<=1;bcd2<=4;bcd1<=5;bcd0<=9; end
			1460: begin bcd3<=1;bcd2<=4;bcd1<=6;bcd0<=0; end
			1461: begin bcd3<=1;bcd2<=4;bcd1<=6;bcd0<=1; end
			1462: begin bcd3<=1;bcd2<=4;bcd1<=6;bcd0<=2; end
			1463: begin bcd3<=1;bcd2<=4;bcd1<=6;bcd0<=3; end
			1464: begin bcd3<=1;bcd2<=4;bcd1<=6;bcd0<=4; end
			1465: begin bcd3<=1;bcd2<=4;bcd1<=6;bcd0<=5; end
			1466: begin bcd3<=1;bcd2<=4;bcd1<=6;bcd0<=6; end
			1467: begin bcd3<=1;bcd2<=4;bcd1<=6;bcd0<=7; end
			1468: begin bcd3<=1;bcd2<=4;bcd1<=6;bcd0<=8; end
			1469: begin bcd3<=1;bcd2<=4;bcd1<=6;bcd0<=9; end
			1470: begin bcd3<=1;bcd2<=4;bcd1<=7;bcd0<=0; end
			1471: begin bcd3<=1;bcd2<=4;bcd1<=7;bcd0<=1; end
			1472: begin bcd3<=1;bcd2<=4;bcd1<=7;bcd0<=2; end
			1473: begin bcd3<=1;bcd2<=4;bcd1<=7;bcd0<=3; end
			1474: begin bcd3<=1;bcd2<=4;bcd1<=7;bcd0<=4; end
			1475: begin bcd3<=1;bcd2<=4;bcd1<=7;bcd0<=5; end
			1476: begin bcd3<=1;bcd2<=4;bcd1<=7;bcd0<=6; end
			1477: begin bcd3<=1;bcd2<=4;bcd1<=7;bcd0<=7; end
			1478: begin bcd3<=1;bcd2<=4;bcd1<=7;bcd0<=8; end
			1479: begin bcd3<=1;bcd2<=4;bcd1<=7;bcd0<=9; end
			1480: begin bcd3<=1;bcd2<=4;bcd1<=8;bcd0<=0; end
			1481: begin bcd3<=1;bcd2<=4;bcd1<=8;bcd0<=1; end
			1482: begin bcd3<=1;bcd2<=4;bcd1<=8;bcd0<=2; end
			1483: begin bcd3<=1;bcd2<=4;bcd1<=8;bcd0<=3; end
			1484: begin bcd3<=1;bcd2<=4;bcd1<=8;bcd0<=4; end
			1485: begin bcd3<=1;bcd2<=4;bcd1<=8;bcd0<=5; end
			1486: begin bcd3<=1;bcd2<=4;bcd1<=8;bcd0<=6; end
			1487: begin bcd3<=1;bcd2<=4;bcd1<=8;bcd0<=7; end
			1488: begin bcd3<=1;bcd2<=4;bcd1<=8;bcd0<=8; end
			1489: begin bcd3<=1;bcd2<=4;bcd1<=8;bcd0<=9; end
			1490: begin bcd3<=1;bcd2<=4;bcd1<=9;bcd0<=0; end
			1491: begin bcd3<=1;bcd2<=4;bcd1<=9;bcd0<=1; end
			1492: begin bcd3<=1;bcd2<=4;bcd1<=9;bcd0<=2; end
			1493: begin bcd3<=1;bcd2<=4;bcd1<=9;bcd0<=3; end
			1494: begin bcd3<=1;bcd2<=4;bcd1<=9;bcd0<=4; end
			1495: begin bcd3<=1;bcd2<=4;bcd1<=9;bcd0<=5; end
			1496: begin bcd3<=1;bcd2<=4;bcd1<=9;bcd0<=6; end
			1497: begin bcd3<=1;bcd2<=4;bcd1<=9;bcd0<=7; end
			1498: begin bcd3<=1;bcd2<=4;bcd1<=9;bcd0<=8; end
			1499: begin bcd3<=1;bcd2<=4;bcd1<=9;bcd0<=9; end
			1500: begin bcd3<=1;bcd2<=5;bcd1<=0;bcd0<=0; end
			1501: begin bcd3<=1;bcd2<=5;bcd1<=0;bcd0<=1; end
			1502: begin bcd3<=1;bcd2<=5;bcd1<=0;bcd0<=2; end
			1503: begin bcd3<=1;bcd2<=5;bcd1<=0;bcd0<=3; end
			1504: begin bcd3<=1;bcd2<=5;bcd1<=0;bcd0<=4; end
			1505: begin bcd3<=1;bcd2<=5;bcd1<=0;bcd0<=5; end
			1506: begin bcd3<=1;bcd2<=5;bcd1<=0;bcd0<=6; end
			1507: begin bcd3<=1;bcd2<=5;bcd1<=0;bcd0<=7; end
			1508: begin bcd3<=1;bcd2<=5;bcd1<=0;bcd0<=8; end
			1509: begin bcd3<=1;bcd2<=5;bcd1<=0;bcd0<=9; end
			1510: begin bcd3<=1;bcd2<=5;bcd1<=1;bcd0<=0; end
			1511: begin bcd3<=1;bcd2<=5;bcd1<=1;bcd0<=1; end
			1512: begin bcd3<=1;bcd2<=5;bcd1<=1;bcd0<=2; end
			1513: begin bcd3<=1;bcd2<=5;bcd1<=1;bcd0<=3; end
			1514: begin bcd3<=1;bcd2<=5;bcd1<=1;bcd0<=4; end
			1515: begin bcd3<=1;bcd2<=5;bcd1<=1;bcd0<=5; end
			1516: begin bcd3<=1;bcd2<=5;bcd1<=1;bcd0<=6; end
			1517: begin bcd3<=1;bcd2<=5;bcd1<=1;bcd0<=7; end
			1518: begin bcd3<=1;bcd2<=5;bcd1<=1;bcd0<=8; end
			1519: begin bcd3<=1;bcd2<=5;bcd1<=1;bcd0<=9; end
			1520: begin bcd3<=1;bcd2<=5;bcd1<=2;bcd0<=0; end
			1521: begin bcd3<=1;bcd2<=5;bcd1<=2;bcd0<=1; end
			1522: begin bcd3<=1;bcd2<=5;bcd1<=2;bcd0<=2; end
			1523: begin bcd3<=1;bcd2<=5;bcd1<=2;bcd0<=3; end
			1524: begin bcd3<=1;bcd2<=5;bcd1<=2;bcd0<=4; end
			1525: begin bcd3<=1;bcd2<=5;bcd1<=2;bcd0<=5; end
			1526: begin bcd3<=1;bcd2<=5;bcd1<=2;bcd0<=6; end
			1527: begin bcd3<=1;bcd2<=5;bcd1<=2;bcd0<=7; end
			1528: begin bcd3<=1;bcd2<=5;bcd1<=2;bcd0<=8; end
			1529: begin bcd3<=1;bcd2<=5;bcd1<=2;bcd0<=9; end
			1530: begin bcd3<=1;bcd2<=5;bcd1<=3;bcd0<=0; end
			1531: begin bcd3<=1;bcd2<=5;bcd1<=3;bcd0<=1; end
			1532: begin bcd3<=1;bcd2<=5;bcd1<=3;bcd0<=2; end
			1533: begin bcd3<=1;bcd2<=5;bcd1<=3;bcd0<=3; end
			1534: begin bcd3<=1;bcd2<=5;bcd1<=3;bcd0<=4; end
			1535: begin bcd3<=1;bcd2<=5;bcd1<=3;bcd0<=5; end
			1536: begin bcd3<=1;bcd2<=5;bcd1<=3;bcd0<=6; end
			1537: begin bcd3<=1;bcd2<=5;bcd1<=3;bcd0<=7; end
			1538: begin bcd3<=1;bcd2<=5;bcd1<=3;bcd0<=8; end
			1539: begin bcd3<=1;bcd2<=5;bcd1<=3;bcd0<=9; end
			1540: begin bcd3<=1;bcd2<=5;bcd1<=4;bcd0<=0; end
			1541: begin bcd3<=1;bcd2<=5;bcd1<=4;bcd0<=1; end
			1542: begin bcd3<=1;bcd2<=5;bcd1<=4;bcd0<=2; end
			1543: begin bcd3<=1;bcd2<=5;bcd1<=4;bcd0<=3; end
			1544: begin bcd3<=1;bcd2<=5;bcd1<=4;bcd0<=4; end
			1545: begin bcd3<=1;bcd2<=5;bcd1<=4;bcd0<=5; end
			1546: begin bcd3<=1;bcd2<=5;bcd1<=4;bcd0<=6; end
			1547: begin bcd3<=1;bcd2<=5;bcd1<=4;bcd0<=7; end
			1548: begin bcd3<=1;bcd2<=5;bcd1<=4;bcd0<=8; end
			1549: begin bcd3<=1;bcd2<=5;bcd1<=4;bcd0<=9; end
			1550: begin bcd3<=1;bcd2<=5;bcd1<=5;bcd0<=0; end
			1551: begin bcd3<=1;bcd2<=5;bcd1<=5;bcd0<=1; end
			1552: begin bcd3<=1;bcd2<=5;bcd1<=5;bcd0<=2; end
			1553: begin bcd3<=1;bcd2<=5;bcd1<=5;bcd0<=3; end
			1554: begin bcd3<=1;bcd2<=5;bcd1<=5;bcd0<=4; end
			1555: begin bcd3<=1;bcd2<=5;bcd1<=5;bcd0<=5; end
			1556: begin bcd3<=1;bcd2<=5;bcd1<=5;bcd0<=6; end
			1557: begin bcd3<=1;bcd2<=5;bcd1<=5;bcd0<=7; end
			1558: begin bcd3<=1;bcd2<=5;bcd1<=5;bcd0<=8; end
			1559: begin bcd3<=1;bcd2<=5;bcd1<=5;bcd0<=9; end
			1560: begin bcd3<=1;bcd2<=5;bcd1<=6;bcd0<=0; end
			1561: begin bcd3<=1;bcd2<=5;bcd1<=6;bcd0<=1; end
			1562: begin bcd3<=1;bcd2<=5;bcd1<=6;bcd0<=2; end
			1563: begin bcd3<=1;bcd2<=5;bcd1<=6;bcd0<=3; end
			1564: begin bcd3<=1;bcd2<=5;bcd1<=6;bcd0<=4; end
			1565: begin bcd3<=1;bcd2<=5;bcd1<=6;bcd0<=5; end
			1566: begin bcd3<=1;bcd2<=5;bcd1<=6;bcd0<=6; end
			1567: begin bcd3<=1;bcd2<=5;bcd1<=6;bcd0<=7; end
			1568: begin bcd3<=1;bcd2<=5;bcd1<=6;bcd0<=8; end
			1569: begin bcd3<=1;bcd2<=5;bcd1<=6;bcd0<=9; end
			1570: begin bcd3<=1;bcd2<=5;bcd1<=7;bcd0<=0; end
			1571: begin bcd3<=1;bcd2<=5;bcd1<=7;bcd0<=1; end
			1572: begin bcd3<=1;bcd2<=5;bcd1<=7;bcd0<=2; end
			1573: begin bcd3<=1;bcd2<=5;bcd1<=7;bcd0<=3; end
			1574: begin bcd3<=1;bcd2<=5;bcd1<=7;bcd0<=4; end
			1575: begin bcd3<=1;bcd2<=5;bcd1<=7;bcd0<=5; end
			1576: begin bcd3<=1;bcd2<=5;bcd1<=7;bcd0<=6; end
			1577: begin bcd3<=1;bcd2<=5;bcd1<=7;bcd0<=7; end
			1578: begin bcd3<=1;bcd2<=5;bcd1<=7;bcd0<=8; end
			1579: begin bcd3<=1;bcd2<=5;bcd1<=7;bcd0<=9; end
			1580: begin bcd3<=1;bcd2<=5;bcd1<=8;bcd0<=0; end
			1581: begin bcd3<=1;bcd2<=5;bcd1<=8;bcd0<=1; end
			1582: begin bcd3<=1;bcd2<=5;bcd1<=8;bcd0<=2; end
			1583: begin bcd3<=1;bcd2<=5;bcd1<=8;bcd0<=3; end
			1584: begin bcd3<=1;bcd2<=5;bcd1<=8;bcd0<=4; end
			1585: begin bcd3<=1;bcd2<=5;bcd1<=8;bcd0<=5; end
			1586: begin bcd3<=1;bcd2<=5;bcd1<=8;bcd0<=6; end
			1587: begin bcd3<=1;bcd2<=5;bcd1<=8;bcd0<=7; end
			1588: begin bcd3<=1;bcd2<=5;bcd1<=8;bcd0<=8; end
			1589: begin bcd3<=1;bcd2<=5;bcd1<=8;bcd0<=9; end
			1590: begin bcd3<=1;bcd2<=5;bcd1<=9;bcd0<=0; end
			1591: begin bcd3<=1;bcd2<=5;bcd1<=9;bcd0<=1; end
			1592: begin bcd3<=1;bcd2<=5;bcd1<=9;bcd0<=2; end
			1593: begin bcd3<=1;bcd2<=5;bcd1<=9;bcd0<=3; end
			1594: begin bcd3<=1;bcd2<=5;bcd1<=9;bcd0<=4; end
			1595: begin bcd3<=1;bcd2<=5;bcd1<=9;bcd0<=5; end
			1596: begin bcd3<=1;bcd2<=5;bcd1<=9;bcd0<=6; end
			1597: begin bcd3<=1;bcd2<=5;bcd1<=9;bcd0<=7; end
			1598: begin bcd3<=1;bcd2<=5;bcd1<=9;bcd0<=8; end
			1599: begin bcd3<=1;bcd2<=5;bcd1<=9;bcd0<=9; end
			1600: begin bcd3<=1;bcd2<=6;bcd1<=0;bcd0<=0; end
			1601: begin bcd3<=1;bcd2<=6;bcd1<=0;bcd0<=1; end
			1602: begin bcd3<=1;bcd2<=6;bcd1<=0;bcd0<=2; end
			1603: begin bcd3<=1;bcd2<=6;bcd1<=0;bcd0<=3; end
			1604: begin bcd3<=1;bcd2<=6;bcd1<=0;bcd0<=4; end
			1605: begin bcd3<=1;bcd2<=6;bcd1<=0;bcd0<=5; end
			1606: begin bcd3<=1;bcd2<=6;bcd1<=0;bcd0<=6; end
			1607: begin bcd3<=1;bcd2<=6;bcd1<=0;bcd0<=7; end
			1608: begin bcd3<=1;bcd2<=6;bcd1<=0;bcd0<=8; end
			1609: begin bcd3<=1;bcd2<=6;bcd1<=0;bcd0<=9; end
			1610: begin bcd3<=1;bcd2<=6;bcd1<=1;bcd0<=0; end
			1611: begin bcd3<=1;bcd2<=6;bcd1<=1;bcd0<=1; end
			1612: begin bcd3<=1;bcd2<=6;bcd1<=1;bcd0<=2; end
			1613: begin bcd3<=1;bcd2<=6;bcd1<=1;bcd0<=3; end
			1614: begin bcd3<=1;bcd2<=6;bcd1<=1;bcd0<=4; end
			1615: begin bcd3<=1;bcd2<=6;bcd1<=1;bcd0<=5; end
			1616: begin bcd3<=1;bcd2<=6;bcd1<=1;bcd0<=6; end
			1617: begin bcd3<=1;bcd2<=6;bcd1<=1;bcd0<=7; end
			1618: begin bcd3<=1;bcd2<=6;bcd1<=1;bcd0<=8; end
			1619: begin bcd3<=1;bcd2<=6;bcd1<=1;bcd0<=9; end
			1620: begin bcd3<=1;bcd2<=6;bcd1<=2;bcd0<=0; end
			1621: begin bcd3<=1;bcd2<=6;bcd1<=2;bcd0<=1; end
			1622: begin bcd3<=1;bcd2<=6;bcd1<=2;bcd0<=2; end
			1623: begin bcd3<=1;bcd2<=6;bcd1<=2;bcd0<=3; end
			1624: begin bcd3<=1;bcd2<=6;bcd1<=2;bcd0<=4; end
			1625: begin bcd3<=1;bcd2<=6;bcd1<=2;bcd0<=5; end
			1626: begin bcd3<=1;bcd2<=6;bcd1<=2;bcd0<=6; end
			1627: begin bcd3<=1;bcd2<=6;bcd1<=2;bcd0<=7; end
			1628: begin bcd3<=1;bcd2<=6;bcd1<=2;bcd0<=8; end
			1629: begin bcd3<=1;bcd2<=6;bcd1<=2;bcd0<=9; end
			1630: begin bcd3<=1;bcd2<=6;bcd1<=3;bcd0<=0; end
			1631: begin bcd3<=1;bcd2<=6;bcd1<=3;bcd0<=1; end
			1632: begin bcd3<=1;bcd2<=6;bcd1<=3;bcd0<=2; end
			1633: begin bcd3<=1;bcd2<=6;bcd1<=3;bcd0<=3; end
			1634: begin bcd3<=1;bcd2<=6;bcd1<=3;bcd0<=4; end
			1635: begin bcd3<=1;bcd2<=6;bcd1<=3;bcd0<=5; end
			1636: begin bcd3<=1;bcd2<=6;bcd1<=3;bcd0<=6; end
			1637: begin bcd3<=1;bcd2<=6;bcd1<=3;bcd0<=7; end
			1638: begin bcd3<=1;bcd2<=6;bcd1<=3;bcd0<=8; end
			1639: begin bcd3<=1;bcd2<=6;bcd1<=3;bcd0<=9; end
			1640: begin bcd3<=1;bcd2<=6;bcd1<=4;bcd0<=0; end
			1641: begin bcd3<=1;bcd2<=6;bcd1<=4;bcd0<=1; end
			1642: begin bcd3<=1;bcd2<=6;bcd1<=4;bcd0<=2; end
			1643: begin bcd3<=1;bcd2<=6;bcd1<=4;bcd0<=3; end
			1644: begin bcd3<=1;bcd2<=6;bcd1<=4;bcd0<=4; end
			1645: begin bcd3<=1;bcd2<=6;bcd1<=4;bcd0<=5; end
			1646: begin bcd3<=1;bcd2<=6;bcd1<=4;bcd0<=6; end
			1647: begin bcd3<=1;bcd2<=6;bcd1<=4;bcd0<=7; end
			1648: begin bcd3<=1;bcd2<=6;bcd1<=4;bcd0<=8; end
			1649: begin bcd3<=1;bcd2<=6;bcd1<=4;bcd0<=9; end
			1650: begin bcd3<=1;bcd2<=6;bcd1<=5;bcd0<=0; end
			1651: begin bcd3<=1;bcd2<=6;bcd1<=5;bcd0<=1; end
			1652: begin bcd3<=1;bcd2<=6;bcd1<=5;bcd0<=2; end
			1653: begin bcd3<=1;bcd2<=6;bcd1<=5;bcd0<=3; end
			1654: begin bcd3<=1;bcd2<=6;bcd1<=5;bcd0<=4; end
			1655: begin bcd3<=1;bcd2<=6;bcd1<=5;bcd0<=5; end
			1656: begin bcd3<=1;bcd2<=6;bcd1<=5;bcd0<=6; end
			1657: begin bcd3<=1;bcd2<=6;bcd1<=5;bcd0<=7; end
			1658: begin bcd3<=1;bcd2<=6;bcd1<=5;bcd0<=8; end
			1659: begin bcd3<=1;bcd2<=6;bcd1<=5;bcd0<=9; end
			1660: begin bcd3<=1;bcd2<=6;bcd1<=6;bcd0<=0; end
			1661: begin bcd3<=1;bcd2<=6;bcd1<=6;bcd0<=1; end
			1662: begin bcd3<=1;bcd2<=6;bcd1<=6;bcd0<=2; end
			1663: begin bcd3<=1;bcd2<=6;bcd1<=6;bcd0<=3; end
			1664: begin bcd3<=1;bcd2<=6;bcd1<=6;bcd0<=4; end
			1665: begin bcd3<=1;bcd2<=6;bcd1<=6;bcd0<=5; end
			1666: begin bcd3<=1;bcd2<=6;bcd1<=6;bcd0<=6; end
			1667: begin bcd3<=1;bcd2<=6;bcd1<=6;bcd0<=7; end
			1668: begin bcd3<=1;bcd2<=6;bcd1<=6;bcd0<=8; end
			1669: begin bcd3<=1;bcd2<=6;bcd1<=6;bcd0<=9; end
			1670: begin bcd3<=1;bcd2<=6;bcd1<=7;bcd0<=0; end
			1671: begin bcd3<=1;bcd2<=6;bcd1<=7;bcd0<=1; end
			1672: begin bcd3<=1;bcd2<=6;bcd1<=7;bcd0<=2; end
			1673: begin bcd3<=1;bcd2<=6;bcd1<=7;bcd0<=3; end
			1674: begin bcd3<=1;bcd2<=6;bcd1<=7;bcd0<=4; end
			1675: begin bcd3<=1;bcd2<=6;bcd1<=7;bcd0<=5; end
			1676: begin bcd3<=1;bcd2<=6;bcd1<=7;bcd0<=6; end
			1677: begin bcd3<=1;bcd2<=6;bcd1<=7;bcd0<=7; end
			1678: begin bcd3<=1;bcd2<=6;bcd1<=7;bcd0<=8; end
			1679: begin bcd3<=1;bcd2<=6;bcd1<=7;bcd0<=9; end
			1680: begin bcd3<=1;bcd2<=6;bcd1<=8;bcd0<=0; end
			1681: begin bcd3<=1;bcd2<=6;bcd1<=8;bcd0<=1; end
			1682: begin bcd3<=1;bcd2<=6;bcd1<=8;bcd0<=2; end
			1683: begin bcd3<=1;bcd2<=6;bcd1<=8;bcd0<=3; end
			1684: begin bcd3<=1;bcd2<=6;bcd1<=8;bcd0<=4; end
			1685: begin bcd3<=1;bcd2<=6;bcd1<=8;bcd0<=5; end
			1686: begin bcd3<=1;bcd2<=6;bcd1<=8;bcd0<=6; end
			1687: begin bcd3<=1;bcd2<=6;bcd1<=8;bcd0<=7; end
			1688: begin bcd3<=1;bcd2<=6;bcd1<=8;bcd0<=8; end
			1689: begin bcd3<=1;bcd2<=6;bcd1<=8;bcd0<=9; end
			1690: begin bcd3<=1;bcd2<=6;bcd1<=9;bcd0<=0; end
			1691: begin bcd3<=1;bcd2<=6;bcd1<=9;bcd0<=1; end
			1692: begin bcd3<=1;bcd2<=6;bcd1<=9;bcd0<=2; end
			1693: begin bcd3<=1;bcd2<=6;bcd1<=9;bcd0<=3; end
			1694: begin bcd3<=1;bcd2<=6;bcd1<=9;bcd0<=4; end
			1695: begin bcd3<=1;bcd2<=6;bcd1<=9;bcd0<=5; end
			1696: begin bcd3<=1;bcd2<=6;bcd1<=9;bcd0<=6; end
			1697: begin bcd3<=1;bcd2<=6;bcd1<=9;bcd0<=7; end
			1698: begin bcd3<=1;bcd2<=6;bcd1<=9;bcd0<=8; end
			1699: begin bcd3<=1;bcd2<=6;bcd1<=9;bcd0<=9; end
			1700: begin bcd3<=1;bcd2<=7;bcd1<=0;bcd0<=0; end
			1701: begin bcd3<=1;bcd2<=7;bcd1<=0;bcd0<=1; end
			1702: begin bcd3<=1;bcd2<=7;bcd1<=0;bcd0<=2; end
			1703: begin bcd3<=1;bcd2<=7;bcd1<=0;bcd0<=3; end
			1704: begin bcd3<=1;bcd2<=7;bcd1<=0;bcd0<=4; end
			1705: begin bcd3<=1;bcd2<=7;bcd1<=0;bcd0<=5; end
			1706: begin bcd3<=1;bcd2<=7;bcd1<=0;bcd0<=6; end
			1707: begin bcd3<=1;bcd2<=7;bcd1<=0;bcd0<=7; end
			1708: begin bcd3<=1;bcd2<=7;bcd1<=0;bcd0<=8; end
			1709: begin bcd3<=1;bcd2<=7;bcd1<=0;bcd0<=9; end
			1710: begin bcd3<=1;bcd2<=7;bcd1<=1;bcd0<=0; end
			1711: begin bcd3<=1;bcd2<=7;bcd1<=1;bcd0<=1; end
			1712: begin bcd3<=1;bcd2<=7;bcd1<=1;bcd0<=2; end
			1713: begin bcd3<=1;bcd2<=7;bcd1<=1;bcd0<=3; end
			1714: begin bcd3<=1;bcd2<=7;bcd1<=1;bcd0<=4; end
			1715: begin bcd3<=1;bcd2<=7;bcd1<=1;bcd0<=5; end
			1716: begin bcd3<=1;bcd2<=7;bcd1<=1;bcd0<=6; end
			1717: begin bcd3<=1;bcd2<=7;bcd1<=1;bcd0<=7; end
			1718: begin bcd3<=1;bcd2<=7;bcd1<=1;bcd0<=8; end
			1719: begin bcd3<=1;bcd2<=7;bcd1<=1;bcd0<=9; end
			1720: begin bcd3<=1;bcd2<=7;bcd1<=2;bcd0<=0; end
			1721: begin bcd3<=1;bcd2<=7;bcd1<=2;bcd0<=1; end
			1722: begin bcd3<=1;bcd2<=7;bcd1<=2;bcd0<=2; end
			1723: begin bcd3<=1;bcd2<=7;bcd1<=2;bcd0<=3; end
			1724: begin bcd3<=1;bcd2<=7;bcd1<=2;bcd0<=4; end
			1725: begin bcd3<=1;bcd2<=7;bcd1<=2;bcd0<=5; end
			1726: begin bcd3<=1;bcd2<=7;bcd1<=2;bcd0<=6; end
			1727: begin bcd3<=1;bcd2<=7;bcd1<=2;bcd0<=7; end
			1728: begin bcd3<=1;bcd2<=7;bcd1<=2;bcd0<=8; end
			1729: begin bcd3<=1;bcd2<=7;bcd1<=2;bcd0<=9; end
			1730: begin bcd3<=1;bcd2<=7;bcd1<=3;bcd0<=0; end
			1731: begin bcd3<=1;bcd2<=7;bcd1<=3;bcd0<=1; end
			1732: begin bcd3<=1;bcd2<=7;bcd1<=3;bcd0<=2; end
			1733: begin bcd3<=1;bcd2<=7;bcd1<=3;bcd0<=3; end
			1734: begin bcd3<=1;bcd2<=7;bcd1<=3;bcd0<=4; end
			1735: begin bcd3<=1;bcd2<=7;bcd1<=3;bcd0<=5; end
			1736: begin bcd3<=1;bcd2<=7;bcd1<=3;bcd0<=6; end
			1737: begin bcd3<=1;bcd2<=7;bcd1<=3;bcd0<=7; end
			1738: begin bcd3<=1;bcd2<=7;bcd1<=3;bcd0<=8; end
			1739: begin bcd3<=1;bcd2<=7;bcd1<=3;bcd0<=9; end
			1740: begin bcd3<=1;bcd2<=7;bcd1<=4;bcd0<=0; end
			1741: begin bcd3<=1;bcd2<=7;bcd1<=4;bcd0<=1; end
			1742: begin bcd3<=1;bcd2<=7;bcd1<=4;bcd0<=2; end
			1743: begin bcd3<=1;bcd2<=7;bcd1<=4;bcd0<=3; end
			1744: begin bcd3<=1;bcd2<=7;bcd1<=4;bcd0<=4; end
			1745: begin bcd3<=1;bcd2<=7;bcd1<=4;bcd0<=5; end
			1746: begin bcd3<=1;bcd2<=7;bcd1<=4;bcd0<=6; end
			1747: begin bcd3<=1;bcd2<=7;bcd1<=4;bcd0<=7; end
			1748: begin bcd3<=1;bcd2<=7;bcd1<=4;bcd0<=8; end
			1749: begin bcd3<=1;bcd2<=7;bcd1<=4;bcd0<=9; end
			1750: begin bcd3<=1;bcd2<=7;bcd1<=5;bcd0<=0; end
			1751: begin bcd3<=1;bcd2<=7;bcd1<=5;bcd0<=1; end
			1752: begin bcd3<=1;bcd2<=7;bcd1<=5;bcd0<=2; end
			1753: begin bcd3<=1;bcd2<=7;bcd1<=5;bcd0<=3; end
			1754: begin bcd3<=1;bcd2<=7;bcd1<=5;bcd0<=4; end
			1755: begin bcd3<=1;bcd2<=7;bcd1<=5;bcd0<=5; end
			1756: begin bcd3<=1;bcd2<=7;bcd1<=5;bcd0<=6; end
			1757: begin bcd3<=1;bcd2<=7;bcd1<=5;bcd0<=7; end
			1758: begin bcd3<=1;bcd2<=7;bcd1<=5;bcd0<=8; end
			1759: begin bcd3<=1;bcd2<=7;bcd1<=5;bcd0<=9; end
			1760: begin bcd3<=1;bcd2<=7;bcd1<=6;bcd0<=0; end
			1761: begin bcd3<=1;bcd2<=7;bcd1<=6;bcd0<=1; end
			1762: begin bcd3<=1;bcd2<=7;bcd1<=6;bcd0<=2; end
			1763: begin bcd3<=1;bcd2<=7;bcd1<=6;bcd0<=3; end
			1764: begin bcd3<=1;bcd2<=7;bcd1<=6;bcd0<=4; end
			1765: begin bcd3<=1;bcd2<=7;bcd1<=6;bcd0<=5; end
			1766: begin bcd3<=1;bcd2<=7;bcd1<=6;bcd0<=6; end
			1767: begin bcd3<=1;bcd2<=7;bcd1<=6;bcd0<=7; end
			1768: begin bcd3<=1;bcd2<=7;bcd1<=6;bcd0<=8; end
			1769: begin bcd3<=1;bcd2<=7;bcd1<=6;bcd0<=9; end
			1770: begin bcd3<=1;bcd2<=7;bcd1<=7;bcd0<=0; end
			1771: begin bcd3<=1;bcd2<=7;bcd1<=7;bcd0<=1; end
			1772: begin bcd3<=1;bcd2<=7;bcd1<=7;bcd0<=2; end
			1773: begin bcd3<=1;bcd2<=7;bcd1<=7;bcd0<=3; end
			1774: begin bcd3<=1;bcd2<=7;bcd1<=7;bcd0<=4; end
			1775: begin bcd3<=1;bcd2<=7;bcd1<=7;bcd0<=5; end
			1776: begin bcd3<=1;bcd2<=7;bcd1<=7;bcd0<=6; end
			1777: begin bcd3<=1;bcd2<=7;bcd1<=7;bcd0<=7; end
			1778: begin bcd3<=1;bcd2<=7;bcd1<=7;bcd0<=8; end
			1779: begin bcd3<=1;bcd2<=7;bcd1<=7;bcd0<=9; end
			1780: begin bcd3<=1;bcd2<=7;bcd1<=8;bcd0<=0; end
			1781: begin bcd3<=1;bcd2<=7;bcd1<=8;bcd0<=1; end
			1782: begin bcd3<=1;bcd2<=7;bcd1<=8;bcd0<=2; end
			1783: begin bcd3<=1;bcd2<=7;bcd1<=8;bcd0<=3; end
			1784: begin bcd3<=1;bcd2<=7;bcd1<=8;bcd0<=4; end
			1785: begin bcd3<=1;bcd2<=7;bcd1<=8;bcd0<=5; end
			1786: begin bcd3<=1;bcd2<=7;bcd1<=8;bcd0<=6; end
			1787: begin bcd3<=1;bcd2<=7;bcd1<=8;bcd0<=7; end
			1788: begin bcd3<=1;bcd2<=7;bcd1<=8;bcd0<=8; end
			1789: begin bcd3<=1;bcd2<=7;bcd1<=8;bcd0<=9; end
			1790: begin bcd3<=1;bcd2<=7;bcd1<=9;bcd0<=0; end
			1791: begin bcd3<=1;bcd2<=7;bcd1<=9;bcd0<=1; end
			1792: begin bcd3<=1;bcd2<=7;bcd1<=9;bcd0<=2; end
			1793: begin bcd3<=1;bcd2<=7;bcd1<=9;bcd0<=3; end
			1794: begin bcd3<=1;bcd2<=7;bcd1<=9;bcd0<=4; end
			1795: begin bcd3<=1;bcd2<=7;bcd1<=9;bcd0<=5; end
			1796: begin bcd3<=1;bcd2<=7;bcd1<=9;bcd0<=6; end
			1797: begin bcd3<=1;bcd2<=7;bcd1<=9;bcd0<=7; end
			1798: begin bcd3<=1;bcd2<=7;bcd1<=9;bcd0<=8; end
			1799: begin bcd3<=1;bcd2<=7;bcd1<=9;bcd0<=9; end
			1800: begin bcd3<=1;bcd2<=8;bcd1<=0;bcd0<=0; end
			1801: begin bcd3<=1;bcd2<=8;bcd1<=0;bcd0<=1; end
			1802: begin bcd3<=1;bcd2<=8;bcd1<=0;bcd0<=2; end
			1803: begin bcd3<=1;bcd2<=8;bcd1<=0;bcd0<=3; end
			1804: begin bcd3<=1;bcd2<=8;bcd1<=0;bcd0<=4; end
			1805: begin bcd3<=1;bcd2<=8;bcd1<=0;bcd0<=5; end
			1806: begin bcd3<=1;bcd2<=8;bcd1<=0;bcd0<=6; end
			1807: begin bcd3<=1;bcd2<=8;bcd1<=0;bcd0<=7; end
			1808: begin bcd3<=1;bcd2<=8;bcd1<=0;bcd0<=8; end
			1809: begin bcd3<=1;bcd2<=8;bcd1<=0;bcd0<=9; end
			1810: begin bcd3<=1;bcd2<=8;bcd1<=1;bcd0<=0; end
			1811: begin bcd3<=1;bcd2<=8;bcd1<=1;bcd0<=1; end
			1812: begin bcd3<=1;bcd2<=8;bcd1<=1;bcd0<=2; end
			1813: begin bcd3<=1;bcd2<=8;bcd1<=1;bcd0<=3; end
			1814: begin bcd3<=1;bcd2<=8;bcd1<=1;bcd0<=4; end
			1815: begin bcd3<=1;bcd2<=8;bcd1<=1;bcd0<=5; end
			1816: begin bcd3<=1;bcd2<=8;bcd1<=1;bcd0<=6; end
			1817: begin bcd3<=1;bcd2<=8;bcd1<=1;bcd0<=7; end
			1818: begin bcd3<=1;bcd2<=8;bcd1<=1;bcd0<=8; end
			1819: begin bcd3<=1;bcd2<=8;bcd1<=1;bcd0<=9; end
			1820: begin bcd3<=1;bcd2<=8;bcd1<=2;bcd0<=0; end
			1821: begin bcd3<=1;bcd2<=8;bcd1<=2;bcd0<=1; end
			1822: begin bcd3<=1;bcd2<=8;bcd1<=2;bcd0<=2; end
			1823: begin bcd3<=1;bcd2<=8;bcd1<=2;bcd0<=3; end
			1824: begin bcd3<=1;bcd2<=8;bcd1<=2;bcd0<=4; end
			1825: begin bcd3<=1;bcd2<=8;bcd1<=2;bcd0<=5; end
			1826: begin bcd3<=1;bcd2<=8;bcd1<=2;bcd0<=6; end
			1827: begin bcd3<=1;bcd2<=8;bcd1<=2;bcd0<=7; end
			1828: begin bcd3<=1;bcd2<=8;bcd1<=2;bcd0<=8; end
			1829: begin bcd3<=1;bcd2<=8;bcd1<=2;bcd0<=9; end
			1830: begin bcd3<=1;bcd2<=8;bcd1<=3;bcd0<=0; end
			1831: begin bcd3<=1;bcd2<=8;bcd1<=3;bcd0<=1; end
			1832: begin bcd3<=1;bcd2<=8;bcd1<=3;bcd0<=2; end
			1833: begin bcd3<=1;bcd2<=8;bcd1<=3;bcd0<=3; end
			1834: begin bcd3<=1;bcd2<=8;bcd1<=3;bcd0<=4; end
			1835: begin bcd3<=1;bcd2<=8;bcd1<=3;bcd0<=5; end
			1836: begin bcd3<=1;bcd2<=8;bcd1<=3;bcd0<=6; end
			1837: begin bcd3<=1;bcd2<=8;bcd1<=3;bcd0<=7; end
			1838: begin bcd3<=1;bcd2<=8;bcd1<=3;bcd0<=8; end
			1839: begin bcd3<=1;bcd2<=8;bcd1<=3;bcd0<=9; end
			1840: begin bcd3<=1;bcd2<=8;bcd1<=4;bcd0<=0; end
			1841: begin bcd3<=1;bcd2<=8;bcd1<=4;bcd0<=1; end
			1842: begin bcd3<=1;bcd2<=8;bcd1<=4;bcd0<=2; end
			1843: begin bcd3<=1;bcd2<=8;bcd1<=4;bcd0<=3; end
			1844: begin bcd3<=1;bcd2<=8;bcd1<=4;bcd0<=4; end
			1845: begin bcd3<=1;bcd2<=8;bcd1<=4;bcd0<=5; end
			1846: begin bcd3<=1;bcd2<=8;bcd1<=4;bcd0<=6; end
			1847: begin bcd3<=1;bcd2<=8;bcd1<=4;bcd0<=7; end
			1848: begin bcd3<=1;bcd2<=8;bcd1<=4;bcd0<=8; end
			1849: begin bcd3<=1;bcd2<=8;bcd1<=4;bcd0<=9; end
			1850: begin bcd3<=1;bcd2<=8;bcd1<=5;bcd0<=0; end
			1851: begin bcd3<=1;bcd2<=8;bcd1<=5;bcd0<=1; end
			1852: begin bcd3<=1;bcd2<=8;bcd1<=5;bcd0<=2; end
			1853: begin bcd3<=1;bcd2<=8;bcd1<=5;bcd0<=3; end
			1854: begin bcd3<=1;bcd2<=8;bcd1<=5;bcd0<=4; end
			1855: begin bcd3<=1;bcd2<=8;bcd1<=5;bcd0<=5; end
			1856: begin bcd3<=1;bcd2<=8;bcd1<=5;bcd0<=6; end
			1857: begin bcd3<=1;bcd2<=8;bcd1<=5;bcd0<=7; end
			1858: begin bcd3<=1;bcd2<=8;bcd1<=5;bcd0<=8; end
			1859: begin bcd3<=1;bcd2<=8;bcd1<=5;bcd0<=9; end
			1860: begin bcd3<=1;bcd2<=8;bcd1<=6;bcd0<=0; end
			1861: begin bcd3<=1;bcd2<=8;bcd1<=6;bcd0<=1; end
			1862: begin bcd3<=1;bcd2<=8;bcd1<=6;bcd0<=2; end
			1863: begin bcd3<=1;bcd2<=8;bcd1<=6;bcd0<=3; end
			1864: begin bcd3<=1;bcd2<=8;bcd1<=6;bcd0<=4; end
			1865: begin bcd3<=1;bcd2<=8;bcd1<=6;bcd0<=5; end
			1866: begin bcd3<=1;bcd2<=8;bcd1<=6;bcd0<=6; end
			1867: begin bcd3<=1;bcd2<=8;bcd1<=6;bcd0<=7; end
			1868: begin bcd3<=1;bcd2<=8;bcd1<=6;bcd0<=8; end
			1869: begin bcd3<=1;bcd2<=8;bcd1<=6;bcd0<=9; end
			1870: begin bcd3<=1;bcd2<=8;bcd1<=7;bcd0<=0; end
			1871: begin bcd3<=1;bcd2<=8;bcd1<=7;bcd0<=1; end
			1872: begin bcd3<=1;bcd2<=8;bcd1<=7;bcd0<=2; end
			1873: begin bcd3<=1;bcd2<=8;bcd1<=7;bcd0<=3; end
			1874: begin bcd3<=1;bcd2<=8;bcd1<=7;bcd0<=4; end
			1875: begin bcd3<=1;bcd2<=8;bcd1<=7;bcd0<=5; end
			1876: begin bcd3<=1;bcd2<=8;bcd1<=7;bcd0<=6; end
			1877: begin bcd3<=1;bcd2<=8;bcd1<=7;bcd0<=7; end
			1878: begin bcd3<=1;bcd2<=8;bcd1<=7;bcd0<=8; end
			1879: begin bcd3<=1;bcd2<=8;bcd1<=7;bcd0<=9; end
			1880: begin bcd3<=1;bcd2<=8;bcd1<=8;bcd0<=0; end
			1881: begin bcd3<=1;bcd2<=8;bcd1<=8;bcd0<=1; end
			1882: begin bcd3<=1;bcd2<=8;bcd1<=8;bcd0<=2; end
			1883: begin bcd3<=1;bcd2<=8;bcd1<=8;bcd0<=3; end
			1884: begin bcd3<=1;bcd2<=8;bcd1<=8;bcd0<=4; end
			1885: begin bcd3<=1;bcd2<=8;bcd1<=8;bcd0<=5; end
			1886: begin bcd3<=1;bcd2<=8;bcd1<=8;bcd0<=6; end
			1887: begin bcd3<=1;bcd2<=8;bcd1<=8;bcd0<=7; end
			1888: begin bcd3<=1;bcd2<=8;bcd1<=8;bcd0<=8; end
			1889: begin bcd3<=1;bcd2<=8;bcd1<=8;bcd0<=9; end
			1890: begin bcd3<=1;bcd2<=8;bcd1<=9;bcd0<=0; end
			1891: begin bcd3<=1;bcd2<=8;bcd1<=9;bcd0<=1; end
			1892: begin bcd3<=1;bcd2<=8;bcd1<=9;bcd0<=2; end
			1893: begin bcd3<=1;bcd2<=8;bcd1<=9;bcd0<=3; end
			1894: begin bcd3<=1;bcd2<=8;bcd1<=9;bcd0<=4; end
			1895: begin bcd3<=1;bcd2<=8;bcd1<=9;bcd0<=5; end
			1896: begin bcd3<=1;bcd2<=8;bcd1<=9;bcd0<=6; end
			1897: begin bcd3<=1;bcd2<=8;bcd1<=9;bcd0<=7; end
			1898: begin bcd3<=1;bcd2<=8;bcd1<=9;bcd0<=8; end
			1899: begin bcd3<=1;bcd2<=8;bcd1<=9;bcd0<=9; end
			1900: begin bcd3<=1;bcd2<=9;bcd1<=0;bcd0<=0; end
			1901: begin bcd3<=1;bcd2<=9;bcd1<=0;bcd0<=1; end
			1902: begin bcd3<=1;bcd2<=9;bcd1<=0;bcd0<=2; end
			1903: begin bcd3<=1;bcd2<=9;bcd1<=0;bcd0<=3; end
			1904: begin bcd3<=1;bcd2<=9;bcd1<=0;bcd0<=4; end
			1905: begin bcd3<=1;bcd2<=9;bcd1<=0;bcd0<=5; end
			1906: begin bcd3<=1;bcd2<=9;bcd1<=0;bcd0<=6; end
			1907: begin bcd3<=1;bcd2<=9;bcd1<=0;bcd0<=7; end
			1908: begin bcd3<=1;bcd2<=9;bcd1<=0;bcd0<=8; end
			1909: begin bcd3<=1;bcd2<=9;bcd1<=0;bcd0<=9; end
			1910: begin bcd3<=1;bcd2<=9;bcd1<=1;bcd0<=0; end
			1911: begin bcd3<=1;bcd2<=9;bcd1<=1;bcd0<=1; end
			1912: begin bcd3<=1;bcd2<=9;bcd1<=1;bcd0<=2; end
			1913: begin bcd3<=1;bcd2<=9;bcd1<=1;bcd0<=3; end
			1914: begin bcd3<=1;bcd2<=9;bcd1<=1;bcd0<=4; end
			1915: begin bcd3<=1;bcd2<=9;bcd1<=1;bcd0<=5; end
			1916: begin bcd3<=1;bcd2<=9;bcd1<=1;bcd0<=6; end
			1917: begin bcd3<=1;bcd2<=9;bcd1<=1;bcd0<=7; end
			1918: begin bcd3<=1;bcd2<=9;bcd1<=1;bcd0<=8; end
			1919: begin bcd3<=1;bcd2<=9;bcd1<=1;bcd0<=9; end
			1920: begin bcd3<=1;bcd2<=9;bcd1<=2;bcd0<=0; end
			1921: begin bcd3<=1;bcd2<=9;bcd1<=2;bcd0<=1; end
			1922: begin bcd3<=1;bcd2<=9;bcd1<=2;bcd0<=2; end
			1923: begin bcd3<=1;bcd2<=9;bcd1<=2;bcd0<=3; end
			1924: begin bcd3<=1;bcd2<=9;bcd1<=2;bcd0<=4; end
			1925: begin bcd3<=1;bcd2<=9;bcd1<=2;bcd0<=5; end
			1926: begin bcd3<=1;bcd2<=9;bcd1<=2;bcd0<=6; end
			1927: begin bcd3<=1;bcd2<=9;bcd1<=2;bcd0<=7; end
			1928: begin bcd3<=1;bcd2<=9;bcd1<=2;bcd0<=8; end
			1929: begin bcd3<=1;bcd2<=9;bcd1<=2;bcd0<=9; end
			1930: begin bcd3<=1;bcd2<=9;bcd1<=3;bcd0<=0; end
			1931: begin bcd3<=1;bcd2<=9;bcd1<=3;bcd0<=1; end
			1932: begin bcd3<=1;bcd2<=9;bcd1<=3;bcd0<=2; end
			1933: begin bcd3<=1;bcd2<=9;bcd1<=3;bcd0<=3; end
			1934: begin bcd3<=1;bcd2<=9;bcd1<=3;bcd0<=4; end
			1935: begin bcd3<=1;bcd2<=9;bcd1<=3;bcd0<=5; end
			1936: begin bcd3<=1;bcd2<=9;bcd1<=3;bcd0<=6; end
			1937: begin bcd3<=1;bcd2<=9;bcd1<=3;bcd0<=7; end
			1938: begin bcd3<=1;bcd2<=9;bcd1<=3;bcd0<=8; end
			1939: begin bcd3<=1;bcd2<=9;bcd1<=3;bcd0<=9; end
			1940: begin bcd3<=1;bcd2<=9;bcd1<=4;bcd0<=0; end
			1941: begin bcd3<=1;bcd2<=9;bcd1<=4;bcd0<=1; end
			1942: begin bcd3<=1;bcd2<=9;bcd1<=4;bcd0<=2; end
			1943: begin bcd3<=1;bcd2<=9;bcd1<=4;bcd0<=3; end
			1944: begin bcd3<=1;bcd2<=9;bcd1<=4;bcd0<=4; end
			1945: begin bcd3<=1;bcd2<=9;bcd1<=4;bcd0<=5; end
			1946: begin bcd3<=1;bcd2<=9;bcd1<=4;bcd0<=6; end
			1947: begin bcd3<=1;bcd2<=9;bcd1<=4;bcd0<=7; end
			1948: begin bcd3<=1;bcd2<=9;bcd1<=4;bcd0<=8; end
			1949: begin bcd3<=1;bcd2<=9;bcd1<=4;bcd0<=9; end
			1950: begin bcd3<=1;bcd2<=9;bcd1<=5;bcd0<=0; end
			1951: begin bcd3<=1;bcd2<=9;bcd1<=5;bcd0<=1; end
			1952: begin bcd3<=1;bcd2<=9;bcd1<=5;bcd0<=2; end
			1953: begin bcd3<=1;bcd2<=9;bcd1<=5;bcd0<=3; end
			1954: begin bcd3<=1;bcd2<=9;bcd1<=5;bcd0<=4; end
			1955: begin bcd3<=1;bcd2<=9;bcd1<=5;bcd0<=5; end
			1956: begin bcd3<=1;bcd2<=9;bcd1<=5;bcd0<=6; end
			1957: begin bcd3<=1;bcd2<=9;bcd1<=5;bcd0<=7; end
			1958: begin bcd3<=1;bcd2<=9;bcd1<=5;bcd0<=8; end
			1959: begin bcd3<=1;bcd2<=9;bcd1<=5;bcd0<=9; end
			1960: begin bcd3<=1;bcd2<=9;bcd1<=6;bcd0<=0; end
			1961: begin bcd3<=1;bcd2<=9;bcd1<=6;bcd0<=1; end
			1962: begin bcd3<=1;bcd2<=9;bcd1<=6;bcd0<=2; end
			1963: begin bcd3<=1;bcd2<=9;bcd1<=6;bcd0<=3; end
			1964: begin bcd3<=1;bcd2<=9;bcd1<=6;bcd0<=4; end
			1965: begin bcd3<=1;bcd2<=9;bcd1<=6;bcd0<=5; end
			1966: begin bcd3<=1;bcd2<=9;bcd1<=6;bcd0<=6; end
			1967: begin bcd3<=1;bcd2<=9;bcd1<=6;bcd0<=7; end
			1968: begin bcd3<=1;bcd2<=9;bcd1<=6;bcd0<=8; end
			1969: begin bcd3<=1;bcd2<=9;bcd1<=6;bcd0<=9; end
			1970: begin bcd3<=1;bcd2<=9;bcd1<=7;bcd0<=0; end
			1971: begin bcd3<=1;bcd2<=9;bcd1<=7;bcd0<=1; end
			1972: begin bcd3<=1;bcd2<=9;bcd1<=7;bcd0<=2; end
			1973: begin bcd3<=1;bcd2<=9;bcd1<=7;bcd0<=3; end
			1974: begin bcd3<=1;bcd2<=9;bcd1<=7;bcd0<=4; end
			1975: begin bcd3<=1;bcd2<=9;bcd1<=7;bcd0<=5; end
			1976: begin bcd3<=1;bcd2<=9;bcd1<=7;bcd0<=6; end
			1977: begin bcd3<=1;bcd2<=9;bcd1<=7;bcd0<=7; end
			1978: begin bcd3<=1;bcd2<=9;bcd1<=7;bcd0<=8; end
			1979: begin bcd3<=1;bcd2<=9;bcd1<=7;bcd0<=9; end
			1980: begin bcd3<=1;bcd2<=9;bcd1<=8;bcd0<=0; end
			1981: begin bcd3<=1;bcd2<=9;bcd1<=8;bcd0<=1; end
			1982: begin bcd3<=1;bcd2<=9;bcd1<=8;bcd0<=2; end
			1983: begin bcd3<=1;bcd2<=9;bcd1<=8;bcd0<=3; end
			1984: begin bcd3<=1;bcd2<=9;bcd1<=8;bcd0<=4; end
			1985: begin bcd3<=1;bcd2<=9;bcd1<=8;bcd0<=5; end
			1986: begin bcd3<=1;bcd2<=9;bcd1<=8;bcd0<=6; end
			1987: begin bcd3<=1;bcd2<=9;bcd1<=8;bcd0<=7; end
			1988: begin bcd3<=1;bcd2<=9;bcd1<=8;bcd0<=8; end
			1989: begin bcd3<=1;bcd2<=9;bcd1<=8;bcd0<=9; end
			1990: begin bcd3<=1;bcd2<=9;bcd1<=9;bcd0<=0; end
			1991: begin bcd3<=1;bcd2<=9;bcd1<=9;bcd0<=1; end
			1992: begin bcd3<=1;bcd2<=9;bcd1<=9;bcd0<=2; end
			1993: begin bcd3<=1;bcd2<=9;bcd1<=9;bcd0<=3; end
			1994: begin bcd3<=1;bcd2<=9;bcd1<=9;bcd0<=4; end
			1995: begin bcd3<=1;bcd2<=9;bcd1<=9;bcd0<=5; end
			1996: begin bcd3<=1;bcd2<=9;bcd1<=9;bcd0<=6; end
			1997: begin bcd3<=1;bcd2<=9;bcd1<=9;bcd0<=7; end
			1998: begin bcd3<=1;bcd2<=9;bcd1<=9;bcd0<=8; end
			1999: begin bcd3<=1;bcd2<=9;bcd1<=9;bcd0<=9; end
			2000: begin bcd3<=2;bcd2<=0;bcd1<=0;bcd0<=0; end
			2001: begin bcd3<=2;bcd2<=0;bcd1<=0;bcd0<=1; end
			2002: begin bcd3<=2;bcd2<=0;bcd1<=0;bcd0<=2; end
			2003: begin bcd3<=2;bcd2<=0;bcd1<=0;bcd0<=3; end
			2004: begin bcd3<=2;bcd2<=0;bcd1<=0;bcd0<=4; end
			2005: begin bcd3<=2;bcd2<=0;bcd1<=0;bcd0<=5; end
			2006: begin bcd3<=2;bcd2<=0;bcd1<=0;bcd0<=6; end
			2007: begin bcd3<=2;bcd2<=0;bcd1<=0;bcd0<=7; end
			2008: begin bcd3<=2;bcd2<=0;bcd1<=0;bcd0<=8; end
			2009: begin bcd3<=2;bcd2<=0;bcd1<=0;bcd0<=9; end
			2010: begin bcd3<=2;bcd2<=0;bcd1<=1;bcd0<=0; end
			2011: begin bcd3<=2;bcd2<=0;bcd1<=1;bcd0<=1; end
			2012: begin bcd3<=2;bcd2<=0;bcd1<=1;bcd0<=2; end
			2013: begin bcd3<=2;bcd2<=0;bcd1<=1;bcd0<=3; end
			2014: begin bcd3<=2;bcd2<=0;bcd1<=1;bcd0<=4; end
			2015: begin bcd3<=2;bcd2<=0;bcd1<=1;bcd0<=5; end
			2016: begin bcd3<=2;bcd2<=0;bcd1<=1;bcd0<=6; end
			2017: begin bcd3<=2;bcd2<=0;bcd1<=1;bcd0<=7; end
			2018: begin bcd3<=2;bcd2<=0;bcd1<=1;bcd0<=8; end
			2019: begin bcd3<=2;bcd2<=0;bcd1<=1;bcd0<=9; end
			2020: begin bcd3<=2;bcd2<=0;bcd1<=2;bcd0<=0; end
			2021: begin bcd3<=2;bcd2<=0;bcd1<=2;bcd0<=1; end
			2022: begin bcd3<=2;bcd2<=0;bcd1<=2;bcd0<=2; end
			2023: begin bcd3<=2;bcd2<=0;bcd1<=2;bcd0<=3; end
			2024: begin bcd3<=2;bcd2<=0;bcd1<=2;bcd0<=4; end
			2025: begin bcd3<=2;bcd2<=0;bcd1<=2;bcd0<=5; end
			2026: begin bcd3<=2;bcd2<=0;bcd1<=2;bcd0<=6; end
			2027: begin bcd3<=2;bcd2<=0;bcd1<=2;bcd0<=7; end
			2028: begin bcd3<=2;bcd2<=0;bcd1<=2;bcd0<=8; end
			2029: begin bcd3<=2;bcd2<=0;bcd1<=2;bcd0<=9; end
			2030: begin bcd3<=2;bcd2<=0;bcd1<=3;bcd0<=0; end
			2031: begin bcd3<=2;bcd2<=0;bcd1<=3;bcd0<=1; end
			2032: begin bcd3<=2;bcd2<=0;bcd1<=3;bcd0<=2; end
			2033: begin bcd3<=2;bcd2<=0;bcd1<=3;bcd0<=3; end
			2034: begin bcd3<=2;bcd2<=0;bcd1<=3;bcd0<=4; end
			2035: begin bcd3<=2;bcd2<=0;bcd1<=3;bcd0<=5; end
			2036: begin bcd3<=2;bcd2<=0;bcd1<=3;bcd0<=6; end
			2037: begin bcd3<=2;bcd2<=0;bcd1<=3;bcd0<=7; end
			2038: begin bcd3<=2;bcd2<=0;bcd1<=3;bcd0<=8; end
			2039: begin bcd3<=2;bcd2<=0;bcd1<=3;bcd0<=9; end
			2040: begin bcd3<=2;bcd2<=0;bcd1<=4;bcd0<=0; end
			2041: begin bcd3<=2;bcd2<=0;bcd1<=4;bcd0<=1; end
			2042: begin bcd3<=2;bcd2<=0;bcd1<=4;bcd0<=2; end
			2043: begin bcd3<=2;bcd2<=0;bcd1<=4;bcd0<=3; end
			2044: begin bcd3<=2;bcd2<=0;bcd1<=4;bcd0<=4; end
			2045: begin bcd3<=2;bcd2<=0;bcd1<=4;bcd0<=5; end
			2046: begin bcd3<=2;bcd2<=0;bcd1<=4;bcd0<=6; end
			2047: begin bcd3<=2;bcd2<=0;bcd1<=4;bcd0<=7; end
			2048: begin bcd3<=2;bcd2<=0;bcd1<=4;bcd0<=8; end
			2049: begin bcd3<=2;bcd2<=0;bcd1<=4;bcd0<=9; end
			2050: begin bcd3<=2;bcd2<=0;bcd1<=5;bcd0<=0; end
			2051: begin bcd3<=2;bcd2<=0;bcd1<=5;bcd0<=1; end
			2052: begin bcd3<=2;bcd2<=0;bcd1<=5;bcd0<=2; end
			2053: begin bcd3<=2;bcd2<=0;bcd1<=5;bcd0<=3; end
			2054: begin bcd3<=2;bcd2<=0;bcd1<=5;bcd0<=4; end
			2055: begin bcd3<=2;bcd2<=0;bcd1<=5;bcd0<=5; end
			2056: begin bcd3<=2;bcd2<=0;bcd1<=5;bcd0<=6; end
			2057: begin bcd3<=2;bcd2<=0;bcd1<=5;bcd0<=7; end
			2058: begin bcd3<=2;bcd2<=0;bcd1<=5;bcd0<=8; end
			2059: begin bcd3<=2;bcd2<=0;bcd1<=5;bcd0<=9; end
			2060: begin bcd3<=2;bcd2<=0;bcd1<=6;bcd0<=0; end
			2061: begin bcd3<=2;bcd2<=0;bcd1<=6;bcd0<=1; end
			2062: begin bcd3<=2;bcd2<=0;bcd1<=6;bcd0<=2; end
			2063: begin bcd3<=2;bcd2<=0;bcd1<=6;bcd0<=3; end
			2064: begin bcd3<=2;bcd2<=0;bcd1<=6;bcd0<=4; end
			2065: begin bcd3<=2;bcd2<=0;bcd1<=6;bcd0<=5; end
			2066: begin bcd3<=2;bcd2<=0;bcd1<=6;bcd0<=6; end
			2067: begin bcd3<=2;bcd2<=0;bcd1<=6;bcd0<=7; end
			2068: begin bcd3<=2;bcd2<=0;bcd1<=6;bcd0<=8; end
			2069: begin bcd3<=2;bcd2<=0;bcd1<=6;bcd0<=9; end
			2070: begin bcd3<=2;bcd2<=0;bcd1<=7;bcd0<=0; end
			2071: begin bcd3<=2;bcd2<=0;bcd1<=7;bcd0<=1; end
			2072: begin bcd3<=2;bcd2<=0;bcd1<=7;bcd0<=2; end
			2073: begin bcd3<=2;bcd2<=0;bcd1<=7;bcd0<=3; end
			2074: begin bcd3<=2;bcd2<=0;bcd1<=7;bcd0<=4; end
			2075: begin bcd3<=2;bcd2<=0;bcd1<=7;bcd0<=5; end
			2076: begin bcd3<=2;bcd2<=0;bcd1<=7;bcd0<=6; end
			2077: begin bcd3<=2;bcd2<=0;bcd1<=7;bcd0<=7; end
			2078: begin bcd3<=2;bcd2<=0;bcd1<=7;bcd0<=8; end
			2079: begin bcd3<=2;bcd2<=0;bcd1<=7;bcd0<=9; end
			2080: begin bcd3<=2;bcd2<=0;bcd1<=8;bcd0<=0; end
			2081: begin bcd3<=2;bcd2<=0;bcd1<=8;bcd0<=1; end
			2082: begin bcd3<=2;bcd2<=0;bcd1<=8;bcd0<=2; end
			2083: begin bcd3<=2;bcd2<=0;bcd1<=8;bcd0<=3; end
			2084: begin bcd3<=2;bcd2<=0;bcd1<=8;bcd0<=4; end
			2085: begin bcd3<=2;bcd2<=0;bcd1<=8;bcd0<=5; end
			2086: begin bcd3<=2;bcd2<=0;bcd1<=8;bcd0<=6; end
			2087: begin bcd3<=2;bcd2<=0;bcd1<=8;bcd0<=7; end
			2088: begin bcd3<=2;bcd2<=0;bcd1<=8;bcd0<=8; end
			2089: begin bcd3<=2;bcd2<=0;bcd1<=8;bcd0<=9; end
			2090: begin bcd3<=2;bcd2<=0;bcd1<=9;bcd0<=0; end
			2091: begin bcd3<=2;bcd2<=0;bcd1<=9;bcd0<=1; end
			2092: begin bcd3<=2;bcd2<=0;bcd1<=9;bcd0<=2; end
			2093: begin bcd3<=2;bcd2<=0;bcd1<=9;bcd0<=3; end
			2094: begin bcd3<=2;bcd2<=0;bcd1<=9;bcd0<=4; end
			2095: begin bcd3<=2;bcd2<=0;bcd1<=9;bcd0<=5; end
			2096: begin bcd3<=2;bcd2<=0;bcd1<=9;bcd0<=6; end
			2097: begin bcd3<=2;bcd2<=0;bcd1<=9;bcd0<=7; end
			2098: begin bcd3<=2;bcd2<=0;bcd1<=9;bcd0<=8; end
			2099: begin bcd3<=2;bcd2<=0;bcd1<=9;bcd0<=9; end
			2100: begin bcd3<=2;bcd2<=1;bcd1<=0;bcd0<=0; end
			2101: begin bcd3<=2;bcd2<=1;bcd1<=0;bcd0<=1; end
			2102: begin bcd3<=2;bcd2<=1;bcd1<=0;bcd0<=2; end
			2103: begin bcd3<=2;bcd2<=1;bcd1<=0;bcd0<=3; end
			2104: begin bcd3<=2;bcd2<=1;bcd1<=0;bcd0<=4; end
			2105: begin bcd3<=2;bcd2<=1;bcd1<=0;bcd0<=5; end
			2106: begin bcd3<=2;bcd2<=1;bcd1<=0;bcd0<=6; end
			2107: begin bcd3<=2;bcd2<=1;bcd1<=0;bcd0<=7; end
			2108: begin bcd3<=2;bcd2<=1;bcd1<=0;bcd0<=8; end
			2109: begin bcd3<=2;bcd2<=1;bcd1<=0;bcd0<=9; end
			2110: begin bcd3<=2;bcd2<=1;bcd1<=1;bcd0<=0; end
			2111: begin bcd3<=2;bcd2<=1;bcd1<=1;bcd0<=1; end
			2112: begin bcd3<=2;bcd2<=1;bcd1<=1;bcd0<=2; end
			2113: begin bcd3<=2;bcd2<=1;bcd1<=1;bcd0<=3; end
			2114: begin bcd3<=2;bcd2<=1;bcd1<=1;bcd0<=4; end
			2115: begin bcd3<=2;bcd2<=1;bcd1<=1;bcd0<=5; end
			2116: begin bcd3<=2;bcd2<=1;bcd1<=1;bcd0<=6; end
			2117: begin bcd3<=2;bcd2<=1;bcd1<=1;bcd0<=7; end
			2118: begin bcd3<=2;bcd2<=1;bcd1<=1;bcd0<=8; end
			2119: begin bcd3<=2;bcd2<=1;bcd1<=1;bcd0<=9; end
			2120: begin bcd3<=2;bcd2<=1;bcd1<=2;bcd0<=0; end
			2121: begin bcd3<=2;bcd2<=1;bcd1<=2;bcd0<=1; end
			2122: begin bcd3<=2;bcd2<=1;bcd1<=2;bcd0<=2; end
			2123: begin bcd3<=2;bcd2<=1;bcd1<=2;bcd0<=3; end
			2124: begin bcd3<=2;bcd2<=1;bcd1<=2;bcd0<=4; end
			2125: begin bcd3<=2;bcd2<=1;bcd1<=2;bcd0<=5; end
			2126: begin bcd3<=2;bcd2<=1;bcd1<=2;bcd0<=6; end
			2127: begin bcd3<=2;bcd2<=1;bcd1<=2;bcd0<=7; end
			2128: begin bcd3<=2;bcd2<=1;bcd1<=2;bcd0<=8; end
			2129: begin bcd3<=2;bcd2<=1;bcd1<=2;bcd0<=9; end
			2130: begin bcd3<=2;bcd2<=1;bcd1<=3;bcd0<=0; end
			2131: begin bcd3<=2;bcd2<=1;bcd1<=3;bcd0<=1; end
			2132: begin bcd3<=2;bcd2<=1;bcd1<=3;bcd0<=2; end
			2133: begin bcd3<=2;bcd2<=1;bcd1<=3;bcd0<=3; end
			2134: begin bcd3<=2;bcd2<=1;bcd1<=3;bcd0<=4; end
			2135: begin bcd3<=2;bcd2<=1;bcd1<=3;bcd0<=5; end
			2136: begin bcd3<=2;bcd2<=1;bcd1<=3;bcd0<=6; end
			2137: begin bcd3<=2;bcd2<=1;bcd1<=3;bcd0<=7; end
			2138: begin bcd3<=2;bcd2<=1;bcd1<=3;bcd0<=8; end
			2139: begin bcd3<=2;bcd2<=1;bcd1<=3;bcd0<=9; end
			2140: begin bcd3<=2;bcd2<=1;bcd1<=4;bcd0<=0; end
			2141: begin bcd3<=2;bcd2<=1;bcd1<=4;bcd0<=1; end
			2142: begin bcd3<=2;bcd2<=1;bcd1<=4;bcd0<=2; end
			2143: begin bcd3<=2;bcd2<=1;bcd1<=4;bcd0<=3; end
			2144: begin bcd3<=2;bcd2<=1;bcd1<=4;bcd0<=4; end
			2145: begin bcd3<=2;bcd2<=1;bcd1<=4;bcd0<=5; end
			2146: begin bcd3<=2;bcd2<=1;bcd1<=4;bcd0<=6; end
			2147: begin bcd3<=2;bcd2<=1;bcd1<=4;bcd0<=7; end
			2148: begin bcd3<=2;bcd2<=1;bcd1<=4;bcd0<=8; end
			2149: begin bcd3<=2;bcd2<=1;bcd1<=4;bcd0<=9; end
			2150: begin bcd3<=2;bcd2<=1;bcd1<=5;bcd0<=0; end
			2151: begin bcd3<=2;bcd2<=1;bcd1<=5;bcd0<=1; end
			2152: begin bcd3<=2;bcd2<=1;bcd1<=5;bcd0<=2; end
			2153: begin bcd3<=2;bcd2<=1;bcd1<=5;bcd0<=3; end
			2154: begin bcd3<=2;bcd2<=1;bcd1<=5;bcd0<=4; end
			2155: begin bcd3<=2;bcd2<=1;bcd1<=5;bcd0<=5; end
			2156: begin bcd3<=2;bcd2<=1;bcd1<=5;bcd0<=6; end
			2157: begin bcd3<=2;bcd2<=1;bcd1<=5;bcd0<=7; end
			2158: begin bcd3<=2;bcd2<=1;bcd1<=5;bcd0<=8; end
			2159: begin bcd3<=2;bcd2<=1;bcd1<=5;bcd0<=9; end
			2160: begin bcd3<=2;bcd2<=1;bcd1<=6;bcd0<=0; end
			2161: begin bcd3<=2;bcd2<=1;bcd1<=6;bcd0<=1; end
			2162: begin bcd3<=2;bcd2<=1;bcd1<=6;bcd0<=2; end
			2163: begin bcd3<=2;bcd2<=1;bcd1<=6;bcd0<=3; end
			2164: begin bcd3<=2;bcd2<=1;bcd1<=6;bcd0<=4; end
			2165: begin bcd3<=2;bcd2<=1;bcd1<=6;bcd0<=5; end
			2166: begin bcd3<=2;bcd2<=1;bcd1<=6;bcd0<=6; end
			2167: begin bcd3<=2;bcd2<=1;bcd1<=6;bcd0<=7; end
			2168: begin bcd3<=2;bcd2<=1;bcd1<=6;bcd0<=8; end
			2169: begin bcd3<=2;bcd2<=1;bcd1<=6;bcd0<=9; end
			2170: begin bcd3<=2;bcd2<=1;bcd1<=7;bcd0<=0; end
			2171: begin bcd3<=2;bcd2<=1;bcd1<=7;bcd0<=1; end
			2172: begin bcd3<=2;bcd2<=1;bcd1<=7;bcd0<=2; end
			2173: begin bcd3<=2;bcd2<=1;bcd1<=7;bcd0<=3; end
			2174: begin bcd3<=2;bcd2<=1;bcd1<=7;bcd0<=4; end
			2175: begin bcd3<=2;bcd2<=1;bcd1<=7;bcd0<=5; end
			2176: begin bcd3<=2;bcd2<=1;bcd1<=7;bcd0<=6; end
			2177: begin bcd3<=2;bcd2<=1;bcd1<=7;bcd0<=7; end
			2178: begin bcd3<=2;bcd2<=1;bcd1<=7;bcd0<=8; end
			2179: begin bcd3<=2;bcd2<=1;bcd1<=7;bcd0<=9; end
			2180: begin bcd3<=2;bcd2<=1;bcd1<=8;bcd0<=0; end
			2181: begin bcd3<=2;bcd2<=1;bcd1<=8;bcd0<=1; end
			2182: begin bcd3<=2;bcd2<=1;bcd1<=8;bcd0<=2; end
			2183: begin bcd3<=2;bcd2<=1;bcd1<=8;bcd0<=3; end
			2184: begin bcd3<=2;bcd2<=1;bcd1<=8;bcd0<=4; end
			2185: begin bcd3<=2;bcd2<=1;bcd1<=8;bcd0<=5; end
			2186: begin bcd3<=2;bcd2<=1;bcd1<=8;bcd0<=6; end
			2187: begin bcd3<=2;bcd2<=1;bcd1<=8;bcd0<=7; end
			2188: begin bcd3<=2;bcd2<=1;bcd1<=8;bcd0<=8; end
			2189: begin bcd3<=2;bcd2<=1;bcd1<=8;bcd0<=9; end
			2190: begin bcd3<=2;bcd2<=1;bcd1<=9;bcd0<=0; end
			2191: begin bcd3<=2;bcd2<=1;bcd1<=9;bcd0<=1; end
			2192: begin bcd3<=2;bcd2<=1;bcd1<=9;bcd0<=2; end
			2193: begin bcd3<=2;bcd2<=1;bcd1<=9;bcd0<=3; end
			2194: begin bcd3<=2;bcd2<=1;bcd1<=9;bcd0<=4; end
			2195: begin bcd3<=2;bcd2<=1;bcd1<=9;bcd0<=5; end
			2196: begin bcd3<=2;bcd2<=1;bcd1<=9;bcd0<=6; end
			2197: begin bcd3<=2;bcd2<=1;bcd1<=9;bcd0<=7; end
			2198: begin bcd3<=2;bcd2<=1;bcd1<=9;bcd0<=8; end
			2199: begin bcd3<=2;bcd2<=1;bcd1<=9;bcd0<=9; end
			2200: begin bcd3<=2;bcd2<=2;bcd1<=0;bcd0<=0; end
			2201: begin bcd3<=2;bcd2<=2;bcd1<=0;bcd0<=1; end
			2202: begin bcd3<=2;bcd2<=2;bcd1<=0;bcd0<=2; end
			2203: begin bcd3<=2;bcd2<=2;bcd1<=0;bcd0<=3; end
			2204: begin bcd3<=2;bcd2<=2;bcd1<=0;bcd0<=4; end
			2205: begin bcd3<=2;bcd2<=2;bcd1<=0;bcd0<=5; end
			2206: begin bcd3<=2;bcd2<=2;bcd1<=0;bcd0<=6; end
			2207: begin bcd3<=2;bcd2<=2;bcd1<=0;bcd0<=7; end
			2208: begin bcd3<=2;bcd2<=2;bcd1<=0;bcd0<=8; end
			2209: begin bcd3<=2;bcd2<=2;bcd1<=0;bcd0<=9; end
			2210: begin bcd3<=2;bcd2<=2;bcd1<=1;bcd0<=0; end
			2211: begin bcd3<=2;bcd2<=2;bcd1<=1;bcd0<=1; end
			2212: begin bcd3<=2;bcd2<=2;bcd1<=1;bcd0<=2; end
			2213: begin bcd3<=2;bcd2<=2;bcd1<=1;bcd0<=3; end
			2214: begin bcd3<=2;bcd2<=2;bcd1<=1;bcd0<=4; end
			2215: begin bcd3<=2;bcd2<=2;bcd1<=1;bcd0<=5; end
			2216: begin bcd3<=2;bcd2<=2;bcd1<=1;bcd0<=6; end
			2217: begin bcd3<=2;bcd2<=2;bcd1<=1;bcd0<=7; end
			2218: begin bcd3<=2;bcd2<=2;bcd1<=1;bcd0<=8; end
			2219: begin bcd3<=2;bcd2<=2;bcd1<=1;bcd0<=9; end
			2220: begin bcd3<=2;bcd2<=2;bcd1<=2;bcd0<=0; end
			2221: begin bcd3<=2;bcd2<=2;bcd1<=2;bcd0<=1; end
			2222: begin bcd3<=2;bcd2<=2;bcd1<=2;bcd0<=2; end
			2223: begin bcd3<=2;bcd2<=2;bcd1<=2;bcd0<=3; end
			2224: begin bcd3<=2;bcd2<=2;bcd1<=2;bcd0<=4; end
			2225: begin bcd3<=2;bcd2<=2;bcd1<=2;bcd0<=5; end
			2226: begin bcd3<=2;bcd2<=2;bcd1<=2;bcd0<=6; end
			2227: begin bcd3<=2;bcd2<=2;bcd1<=2;bcd0<=7; end
			2228: begin bcd3<=2;bcd2<=2;bcd1<=2;bcd0<=8; end
			2229: begin bcd3<=2;bcd2<=2;bcd1<=2;bcd0<=9; end
			2230: begin bcd3<=2;bcd2<=2;bcd1<=3;bcd0<=0; end
			2231: begin bcd3<=2;bcd2<=2;bcd1<=3;bcd0<=1; end
			2232: begin bcd3<=2;bcd2<=2;bcd1<=3;bcd0<=2; end
			2233: begin bcd3<=2;bcd2<=2;bcd1<=3;bcd0<=3; end
			2234: begin bcd3<=2;bcd2<=2;bcd1<=3;bcd0<=4; end
			2235: begin bcd3<=2;bcd2<=2;bcd1<=3;bcd0<=5; end
			2236: begin bcd3<=2;bcd2<=2;bcd1<=3;bcd0<=6; end
			2237: begin bcd3<=2;bcd2<=2;bcd1<=3;bcd0<=7; end
			2238: begin bcd3<=2;bcd2<=2;bcd1<=3;bcd0<=8; end
			2239: begin bcd3<=2;bcd2<=2;bcd1<=3;bcd0<=9; end
			2240: begin bcd3<=2;bcd2<=2;bcd1<=4;bcd0<=0; end
			2241: begin bcd3<=2;bcd2<=2;bcd1<=4;bcd0<=1; end
			2242: begin bcd3<=2;bcd2<=2;bcd1<=4;bcd0<=2; end
			2243: begin bcd3<=2;bcd2<=2;bcd1<=4;bcd0<=3; end
			2244: begin bcd3<=2;bcd2<=2;bcd1<=4;bcd0<=4; end
			2245: begin bcd3<=2;bcd2<=2;bcd1<=4;bcd0<=5; end
			2246: begin bcd3<=2;bcd2<=2;bcd1<=4;bcd0<=6; end
			2247: begin bcd3<=2;bcd2<=2;bcd1<=4;bcd0<=7; end
			2248: begin bcd3<=2;bcd2<=2;bcd1<=4;bcd0<=8; end
			2249: begin bcd3<=2;bcd2<=2;bcd1<=4;bcd0<=9; end
			2250: begin bcd3<=2;bcd2<=2;bcd1<=5;bcd0<=0; end
			2251: begin bcd3<=2;bcd2<=2;bcd1<=5;bcd0<=1; end
			2252: begin bcd3<=2;bcd2<=2;bcd1<=5;bcd0<=2; end
			2253: begin bcd3<=2;bcd2<=2;bcd1<=5;bcd0<=3; end
			2254: begin bcd3<=2;bcd2<=2;bcd1<=5;bcd0<=4; end
			2255: begin bcd3<=2;bcd2<=2;bcd1<=5;bcd0<=5; end
			2256: begin bcd3<=2;bcd2<=2;bcd1<=5;bcd0<=6; end
			2257: begin bcd3<=2;bcd2<=2;bcd1<=5;bcd0<=7; end
			2258: begin bcd3<=2;bcd2<=2;bcd1<=5;bcd0<=8; end
			2259: begin bcd3<=2;bcd2<=2;bcd1<=5;bcd0<=9; end
			2260: begin bcd3<=2;bcd2<=2;bcd1<=6;bcd0<=0; end
			2261: begin bcd3<=2;bcd2<=2;bcd1<=6;bcd0<=1; end
			2262: begin bcd3<=2;bcd2<=2;bcd1<=6;bcd0<=2; end
			2263: begin bcd3<=2;bcd2<=2;bcd1<=6;bcd0<=3; end
			2264: begin bcd3<=2;bcd2<=2;bcd1<=6;bcd0<=4; end
			2265: begin bcd3<=2;bcd2<=2;bcd1<=6;bcd0<=5; end
			2266: begin bcd3<=2;bcd2<=2;bcd1<=6;bcd0<=6; end
			2267: begin bcd3<=2;bcd2<=2;bcd1<=6;bcd0<=7; end
			2268: begin bcd3<=2;bcd2<=2;bcd1<=6;bcd0<=8; end
			2269: begin bcd3<=2;bcd2<=2;bcd1<=6;bcd0<=9; end
			2270: begin bcd3<=2;bcd2<=2;bcd1<=7;bcd0<=0; end
			2271: begin bcd3<=2;bcd2<=2;bcd1<=7;bcd0<=1; end
			2272: begin bcd3<=2;bcd2<=2;bcd1<=7;bcd0<=2; end
			2273: begin bcd3<=2;bcd2<=2;bcd1<=7;bcd0<=3; end
			2274: begin bcd3<=2;bcd2<=2;bcd1<=7;bcd0<=4; end
			2275: begin bcd3<=2;bcd2<=2;bcd1<=7;bcd0<=5; end
			2276: begin bcd3<=2;bcd2<=2;bcd1<=7;bcd0<=6; end
			2277: begin bcd3<=2;bcd2<=2;bcd1<=7;bcd0<=7; end
			2278: begin bcd3<=2;bcd2<=2;bcd1<=7;bcd0<=8; end
			2279: begin bcd3<=2;bcd2<=2;bcd1<=7;bcd0<=9; end
			2280: begin bcd3<=2;bcd2<=2;bcd1<=8;bcd0<=0; end
			2281: begin bcd3<=2;bcd2<=2;bcd1<=8;bcd0<=1; end
			2282: begin bcd3<=2;bcd2<=2;bcd1<=8;bcd0<=2; end
			2283: begin bcd3<=2;bcd2<=2;bcd1<=8;bcd0<=3; end
			2284: begin bcd3<=2;bcd2<=2;bcd1<=8;bcd0<=4; end
			2285: begin bcd3<=2;bcd2<=2;bcd1<=8;bcd0<=5; end
			2286: begin bcd3<=2;bcd2<=2;bcd1<=8;bcd0<=6; end
			2287: begin bcd3<=2;bcd2<=2;bcd1<=8;bcd0<=7; end
			2288: begin bcd3<=2;bcd2<=2;bcd1<=8;bcd0<=8; end
			2289: begin bcd3<=2;bcd2<=2;bcd1<=8;bcd0<=9; end
			2290: begin bcd3<=2;bcd2<=2;bcd1<=9;bcd0<=0; end
			2291: begin bcd3<=2;bcd2<=2;bcd1<=9;bcd0<=1; end
			2292: begin bcd3<=2;bcd2<=2;bcd1<=9;bcd0<=2; end
			2293: begin bcd3<=2;bcd2<=2;bcd1<=9;bcd0<=3; end
			2294: begin bcd3<=2;bcd2<=2;bcd1<=9;bcd0<=4; end
			2295: begin bcd3<=2;bcd2<=2;bcd1<=9;bcd0<=5; end
			2296: begin bcd3<=2;bcd2<=2;bcd1<=9;bcd0<=6; end
			2297: begin bcd3<=2;bcd2<=2;bcd1<=9;bcd0<=7; end
			2298: begin bcd3<=2;bcd2<=2;bcd1<=9;bcd0<=8; end
			2299: begin bcd3<=2;bcd2<=2;bcd1<=9;bcd0<=9; end
			2300: begin bcd3<=2;bcd2<=3;bcd1<=0;bcd0<=0; end
			2301: begin bcd3<=2;bcd2<=3;bcd1<=0;bcd0<=1; end
			2302: begin bcd3<=2;bcd2<=3;bcd1<=0;bcd0<=2; end
			2303: begin bcd3<=2;bcd2<=3;bcd1<=0;bcd0<=3; end
			2304: begin bcd3<=2;bcd2<=3;bcd1<=0;bcd0<=4; end
			2305: begin bcd3<=2;bcd2<=3;bcd1<=0;bcd0<=5; end
			2306: begin bcd3<=2;bcd2<=3;bcd1<=0;bcd0<=6; end
			2307: begin bcd3<=2;bcd2<=3;bcd1<=0;bcd0<=7; end
			2308: begin bcd3<=2;bcd2<=3;bcd1<=0;bcd0<=8; end
			2309: begin bcd3<=2;bcd2<=3;bcd1<=0;bcd0<=9; end
			2310: begin bcd3<=2;bcd2<=3;bcd1<=1;bcd0<=0; end
			2311: begin bcd3<=2;bcd2<=3;bcd1<=1;bcd0<=1; end
			2312: begin bcd3<=2;bcd2<=3;bcd1<=1;bcd0<=2; end
			2313: begin bcd3<=2;bcd2<=3;bcd1<=1;bcd0<=3; end
			2314: begin bcd3<=2;bcd2<=3;bcd1<=1;bcd0<=4; end
			2315: begin bcd3<=2;bcd2<=3;bcd1<=1;bcd0<=5; end
			2316: begin bcd3<=2;bcd2<=3;bcd1<=1;bcd0<=6; end
			2317: begin bcd3<=2;bcd2<=3;bcd1<=1;bcd0<=7; end
			2318: begin bcd3<=2;bcd2<=3;bcd1<=1;bcd0<=8; end
			2319: begin bcd3<=2;bcd2<=3;bcd1<=1;bcd0<=9; end
			2320: begin bcd3<=2;bcd2<=3;bcd1<=2;bcd0<=0; end
			2321: begin bcd3<=2;bcd2<=3;bcd1<=2;bcd0<=1; end
			2322: begin bcd3<=2;bcd2<=3;bcd1<=2;bcd0<=2; end
			2323: begin bcd3<=2;bcd2<=3;bcd1<=2;bcd0<=3; end
			2324: begin bcd3<=2;bcd2<=3;bcd1<=2;bcd0<=4; end
			2325: begin bcd3<=2;bcd2<=3;bcd1<=2;bcd0<=5; end
			2326: begin bcd3<=2;bcd2<=3;bcd1<=2;bcd0<=6; end
			2327: begin bcd3<=2;bcd2<=3;bcd1<=2;bcd0<=7; end
			2328: begin bcd3<=2;bcd2<=3;bcd1<=2;bcd0<=8; end
			2329: begin bcd3<=2;bcd2<=3;bcd1<=2;bcd0<=9; end
			2330: begin bcd3<=2;bcd2<=3;bcd1<=3;bcd0<=0; end
			2331: begin bcd3<=2;bcd2<=3;bcd1<=3;bcd0<=1; end
			2332: begin bcd3<=2;bcd2<=3;bcd1<=3;bcd0<=2; end
			2333: begin bcd3<=2;bcd2<=3;bcd1<=3;bcd0<=3; end
			2334: begin bcd3<=2;bcd2<=3;bcd1<=3;bcd0<=4; end
			2335: begin bcd3<=2;bcd2<=3;bcd1<=3;bcd0<=5; end
			2336: begin bcd3<=2;bcd2<=3;bcd1<=3;bcd0<=6; end
			2337: begin bcd3<=2;bcd2<=3;bcd1<=3;bcd0<=7; end
			2338: begin bcd3<=2;bcd2<=3;bcd1<=3;bcd0<=8; end
			2339: begin bcd3<=2;bcd2<=3;bcd1<=3;bcd0<=9; end
			2340: begin bcd3<=2;bcd2<=3;bcd1<=4;bcd0<=0; end
			2341: begin bcd3<=2;bcd2<=3;bcd1<=4;bcd0<=1; end
			2342: begin bcd3<=2;bcd2<=3;bcd1<=4;bcd0<=2; end
			2343: begin bcd3<=2;bcd2<=3;bcd1<=4;bcd0<=3; end
			2344: begin bcd3<=2;bcd2<=3;bcd1<=4;bcd0<=4; end
			2345: begin bcd3<=2;bcd2<=3;bcd1<=4;bcd0<=5; end
			2346: begin bcd3<=2;bcd2<=3;bcd1<=4;bcd0<=6; end
			2347: begin bcd3<=2;bcd2<=3;bcd1<=4;bcd0<=7; end
			2348: begin bcd3<=2;bcd2<=3;bcd1<=4;bcd0<=8; end
			2349: begin bcd3<=2;bcd2<=3;bcd1<=4;bcd0<=9; end
			2350: begin bcd3<=2;bcd2<=3;bcd1<=5;bcd0<=0; end
			2351: begin bcd3<=2;bcd2<=3;bcd1<=5;bcd0<=1; end
			2352: begin bcd3<=2;bcd2<=3;bcd1<=5;bcd0<=2; end
			2353: begin bcd3<=2;bcd2<=3;bcd1<=5;bcd0<=3; end
			2354: begin bcd3<=2;bcd2<=3;bcd1<=5;bcd0<=4; end
			2355: begin bcd3<=2;bcd2<=3;bcd1<=5;bcd0<=5; end
			2356: begin bcd3<=2;bcd2<=3;bcd1<=5;bcd0<=6; end
			2357: begin bcd3<=2;bcd2<=3;bcd1<=5;bcd0<=7; end
			2358: begin bcd3<=2;bcd2<=3;bcd1<=5;bcd0<=8; end
			2359: begin bcd3<=2;bcd2<=3;bcd1<=5;bcd0<=9; end
			2360: begin bcd3<=2;bcd2<=3;bcd1<=6;bcd0<=0; end
			2361: begin bcd3<=2;bcd2<=3;bcd1<=6;bcd0<=1; end
			2362: begin bcd3<=2;bcd2<=3;bcd1<=6;bcd0<=2; end
			2363: begin bcd3<=2;bcd2<=3;bcd1<=6;bcd0<=3; end
			2364: begin bcd3<=2;bcd2<=3;bcd1<=6;bcd0<=4; end
			2365: begin bcd3<=2;bcd2<=3;bcd1<=6;bcd0<=5; end
			2366: begin bcd3<=2;bcd2<=3;bcd1<=6;bcd0<=6; end
			2367: begin bcd3<=2;bcd2<=3;bcd1<=6;bcd0<=7; end
			2368: begin bcd3<=2;bcd2<=3;bcd1<=6;bcd0<=8; end
			2369: begin bcd3<=2;bcd2<=3;bcd1<=6;bcd0<=9; end
			2370: begin bcd3<=2;bcd2<=3;bcd1<=7;bcd0<=0; end
			2371: begin bcd3<=2;bcd2<=3;bcd1<=7;bcd0<=1; end
			2372: begin bcd3<=2;bcd2<=3;bcd1<=7;bcd0<=2; end
			2373: begin bcd3<=2;bcd2<=3;bcd1<=7;bcd0<=3; end
			2374: begin bcd3<=2;bcd2<=3;bcd1<=7;bcd0<=4; end
			2375: begin bcd3<=2;bcd2<=3;bcd1<=7;bcd0<=5; end
			2376: begin bcd3<=2;bcd2<=3;bcd1<=7;bcd0<=6; end
			2377: begin bcd3<=2;bcd2<=3;bcd1<=7;bcd0<=7; end
			2378: begin bcd3<=2;bcd2<=3;bcd1<=7;bcd0<=8; end
			2379: begin bcd3<=2;bcd2<=3;bcd1<=7;bcd0<=9; end
			2380: begin bcd3<=2;bcd2<=3;bcd1<=8;bcd0<=0; end
			2381: begin bcd3<=2;bcd2<=3;bcd1<=8;bcd0<=1; end
			2382: begin bcd3<=2;bcd2<=3;bcd1<=8;bcd0<=2; end
			2383: begin bcd3<=2;bcd2<=3;bcd1<=8;bcd0<=3; end
			2384: begin bcd3<=2;bcd2<=3;bcd1<=8;bcd0<=4; end
			2385: begin bcd3<=2;bcd2<=3;bcd1<=8;bcd0<=5; end
			2386: begin bcd3<=2;bcd2<=3;bcd1<=8;bcd0<=6; end
			2387: begin bcd3<=2;bcd2<=3;bcd1<=8;bcd0<=7; end
			2388: begin bcd3<=2;bcd2<=3;bcd1<=8;bcd0<=8; end
			2389: begin bcd3<=2;bcd2<=3;bcd1<=8;bcd0<=9; end
			2390: begin bcd3<=2;bcd2<=3;bcd1<=9;bcd0<=0; end
			2391: begin bcd3<=2;bcd2<=3;bcd1<=9;bcd0<=1; end
			2392: begin bcd3<=2;bcd2<=3;bcd1<=9;bcd0<=2; end
			2393: begin bcd3<=2;bcd2<=3;bcd1<=9;bcd0<=3; end
			2394: begin bcd3<=2;bcd2<=3;bcd1<=9;bcd0<=4; end
			2395: begin bcd3<=2;bcd2<=3;bcd1<=9;bcd0<=5; end
			2396: begin bcd3<=2;bcd2<=3;bcd1<=9;bcd0<=6; end
			2397: begin bcd3<=2;bcd2<=3;bcd1<=9;bcd0<=7; end
			2398: begin bcd3<=2;bcd2<=3;bcd1<=9;bcd0<=8; end
			2399: begin bcd3<=2;bcd2<=3;bcd1<=9;bcd0<=9; end
			2400: begin bcd3<=2;bcd2<=4;bcd1<=0;bcd0<=0; end
			2401: begin bcd3<=2;bcd2<=4;bcd1<=0;bcd0<=1; end
			2402: begin bcd3<=2;bcd2<=4;bcd1<=0;bcd0<=2; end
			2403: begin bcd3<=2;bcd2<=4;bcd1<=0;bcd0<=3; end
			2404: begin bcd3<=2;bcd2<=4;bcd1<=0;bcd0<=4; end
			2405: begin bcd3<=2;bcd2<=4;bcd1<=0;bcd0<=5; end
			2406: begin bcd3<=2;bcd2<=4;bcd1<=0;bcd0<=6; end
			2407: begin bcd3<=2;bcd2<=4;bcd1<=0;bcd0<=7; end
			2408: begin bcd3<=2;bcd2<=4;bcd1<=0;bcd0<=8; end
			2409: begin bcd3<=2;bcd2<=4;bcd1<=0;bcd0<=9; end
			2410: begin bcd3<=2;bcd2<=4;bcd1<=1;bcd0<=0; end
			2411: begin bcd3<=2;bcd2<=4;bcd1<=1;bcd0<=1; end
			2412: begin bcd3<=2;bcd2<=4;bcd1<=1;bcd0<=2; end
			2413: begin bcd3<=2;bcd2<=4;bcd1<=1;bcd0<=3; end
			2414: begin bcd3<=2;bcd2<=4;bcd1<=1;bcd0<=4; end
			2415: begin bcd3<=2;bcd2<=4;bcd1<=1;bcd0<=5; end
			2416: begin bcd3<=2;bcd2<=4;bcd1<=1;bcd0<=6; end
			2417: begin bcd3<=2;bcd2<=4;bcd1<=1;bcd0<=7; end
			2418: begin bcd3<=2;bcd2<=4;bcd1<=1;bcd0<=8; end
			2419: begin bcd3<=2;bcd2<=4;bcd1<=1;bcd0<=9; end
			2420: begin bcd3<=2;bcd2<=4;bcd1<=2;bcd0<=0; end
			2421: begin bcd3<=2;bcd2<=4;bcd1<=2;bcd0<=1; end
			2422: begin bcd3<=2;bcd2<=4;bcd1<=2;bcd0<=2; end
			2423: begin bcd3<=2;bcd2<=4;bcd1<=2;bcd0<=3; end
			2424: begin bcd3<=2;bcd2<=4;bcd1<=2;bcd0<=4; end
			2425: begin bcd3<=2;bcd2<=4;bcd1<=2;bcd0<=5; end
			2426: begin bcd3<=2;bcd2<=4;bcd1<=2;bcd0<=6; end
			2427: begin bcd3<=2;bcd2<=4;bcd1<=2;bcd0<=7; end
			2428: begin bcd3<=2;bcd2<=4;bcd1<=2;bcd0<=8; end
			2429: begin bcd3<=2;bcd2<=4;bcd1<=2;bcd0<=9; end
			2430: begin bcd3<=2;bcd2<=4;bcd1<=3;bcd0<=0; end
			2431: begin bcd3<=2;bcd2<=4;bcd1<=3;bcd0<=1; end
			2432: begin bcd3<=2;bcd2<=4;bcd1<=3;bcd0<=2; end
			2433: begin bcd3<=2;bcd2<=4;bcd1<=3;bcd0<=3; end
			2434: begin bcd3<=2;bcd2<=4;bcd1<=3;bcd0<=4; end
			2435: begin bcd3<=2;bcd2<=4;bcd1<=3;bcd0<=5; end
			2436: begin bcd3<=2;bcd2<=4;bcd1<=3;bcd0<=6; end
			2437: begin bcd3<=2;bcd2<=4;bcd1<=3;bcd0<=7; end
			2438: begin bcd3<=2;bcd2<=4;bcd1<=3;bcd0<=8; end
			2439: begin bcd3<=2;bcd2<=4;bcd1<=3;bcd0<=9; end
			2440: begin bcd3<=2;bcd2<=4;bcd1<=4;bcd0<=0; end
			2441: begin bcd3<=2;bcd2<=4;bcd1<=4;bcd0<=1; end
			2442: begin bcd3<=2;bcd2<=4;bcd1<=4;bcd0<=2; end
			2443: begin bcd3<=2;bcd2<=4;bcd1<=4;bcd0<=3; end
			2444: begin bcd3<=2;bcd2<=4;bcd1<=4;bcd0<=4; end
			2445: begin bcd3<=2;bcd2<=4;bcd1<=4;bcd0<=5; end
			2446: begin bcd3<=2;bcd2<=4;bcd1<=4;bcd0<=6; end
			2447: begin bcd3<=2;bcd2<=4;bcd1<=4;bcd0<=7; end
			2448: begin bcd3<=2;bcd2<=4;bcd1<=4;bcd0<=8; end
			2449: begin bcd3<=2;bcd2<=4;bcd1<=4;bcd0<=9; end
			2450: begin bcd3<=2;bcd2<=4;bcd1<=5;bcd0<=0; end
			2451: begin bcd3<=2;bcd2<=4;bcd1<=5;bcd0<=1; end
			2452: begin bcd3<=2;bcd2<=4;bcd1<=5;bcd0<=2; end
			2453: begin bcd3<=2;bcd2<=4;bcd1<=5;bcd0<=3; end
			2454: begin bcd3<=2;bcd2<=4;bcd1<=5;bcd0<=4; end
			2455: begin bcd3<=2;bcd2<=4;bcd1<=5;bcd0<=5; end
			2456: begin bcd3<=2;bcd2<=4;bcd1<=5;bcd0<=6; end
			2457: begin bcd3<=2;bcd2<=4;bcd1<=5;bcd0<=7; end
			2458: begin bcd3<=2;bcd2<=4;bcd1<=5;bcd0<=8; end
			2459: begin bcd3<=2;bcd2<=4;bcd1<=5;bcd0<=9; end
			2460: begin bcd3<=2;bcd2<=4;bcd1<=6;bcd0<=0; end
			2461: begin bcd3<=2;bcd2<=4;bcd1<=6;bcd0<=1; end
			2462: begin bcd3<=2;bcd2<=4;bcd1<=6;bcd0<=2; end
			2463: begin bcd3<=2;bcd2<=4;bcd1<=6;bcd0<=3; end
			2464: begin bcd3<=2;bcd2<=4;bcd1<=6;bcd0<=4; end
			2465: begin bcd3<=2;bcd2<=4;bcd1<=6;bcd0<=5; end
			2466: begin bcd3<=2;bcd2<=4;bcd1<=6;bcd0<=6; end
			2467: begin bcd3<=2;bcd2<=4;bcd1<=6;bcd0<=7; end
			2468: begin bcd3<=2;bcd2<=4;bcd1<=6;bcd0<=8; end
			2469: begin bcd3<=2;bcd2<=4;bcd1<=6;bcd0<=9; end
			2470: begin bcd3<=2;bcd2<=4;bcd1<=7;bcd0<=0; end
			2471: begin bcd3<=2;bcd2<=4;bcd1<=7;bcd0<=1; end
			2472: begin bcd3<=2;bcd2<=4;bcd1<=7;bcd0<=2; end
			2473: begin bcd3<=2;bcd2<=4;bcd1<=7;bcd0<=3; end
			2474: begin bcd3<=2;bcd2<=4;bcd1<=7;bcd0<=4; end
			2475: begin bcd3<=2;bcd2<=4;bcd1<=7;bcd0<=5; end
			2476: begin bcd3<=2;bcd2<=4;bcd1<=7;bcd0<=6; end
			2477: begin bcd3<=2;bcd2<=4;bcd1<=7;bcd0<=7; end
			2478: begin bcd3<=2;bcd2<=4;bcd1<=7;bcd0<=8; end
			2479: begin bcd3<=2;bcd2<=4;bcd1<=7;bcd0<=9; end
			2480: begin bcd3<=2;bcd2<=4;bcd1<=8;bcd0<=0; end
			2481: begin bcd3<=2;bcd2<=4;bcd1<=8;bcd0<=1; end
			2482: begin bcd3<=2;bcd2<=4;bcd1<=8;bcd0<=2; end
			2483: begin bcd3<=2;bcd2<=4;bcd1<=8;bcd0<=3; end
			2484: begin bcd3<=2;bcd2<=4;bcd1<=8;bcd0<=4; end
			2485: begin bcd3<=2;bcd2<=4;bcd1<=8;bcd0<=5; end
			2486: begin bcd3<=2;bcd2<=4;bcd1<=8;bcd0<=6; end
			2487: begin bcd3<=2;bcd2<=4;bcd1<=8;bcd0<=7; end
			2488: begin bcd3<=2;bcd2<=4;bcd1<=8;bcd0<=8; end
			2489: begin bcd3<=2;bcd2<=4;bcd1<=8;bcd0<=9; end
			2490: begin bcd3<=2;bcd2<=4;bcd1<=9;bcd0<=0; end
			2491: begin bcd3<=2;bcd2<=4;bcd1<=9;bcd0<=1; end
			2492: begin bcd3<=2;bcd2<=4;bcd1<=9;bcd0<=2; end
			2493: begin bcd3<=2;bcd2<=4;bcd1<=9;bcd0<=3; end
			2494: begin bcd3<=2;bcd2<=4;bcd1<=9;bcd0<=4; end
			2495: begin bcd3<=2;bcd2<=4;bcd1<=9;bcd0<=5; end
			2496: begin bcd3<=2;bcd2<=4;bcd1<=9;bcd0<=6; end
			2497: begin bcd3<=2;bcd2<=4;bcd1<=9;bcd0<=7; end
			2498: begin bcd3<=2;bcd2<=4;bcd1<=9;bcd0<=8; end
			2499: begin bcd3<=2;bcd2<=4;bcd1<=9;bcd0<=9; end
			2500: begin bcd3<=2;bcd2<=5;bcd1<=0;bcd0<=0; end
			2501: begin bcd3<=2;bcd2<=5;bcd1<=0;bcd0<=1; end
			2502: begin bcd3<=2;bcd2<=5;bcd1<=0;bcd0<=2; end
			2503: begin bcd3<=2;bcd2<=5;bcd1<=0;bcd0<=3; end
			2504: begin bcd3<=2;bcd2<=5;bcd1<=0;bcd0<=4; end
			2505: begin bcd3<=2;bcd2<=5;bcd1<=0;bcd0<=5; end
			2506: begin bcd3<=2;bcd2<=5;bcd1<=0;bcd0<=6; end
			2507: begin bcd3<=2;bcd2<=5;bcd1<=0;bcd0<=7; end
			2508: begin bcd3<=2;bcd2<=5;bcd1<=0;bcd0<=8; end
			2509: begin bcd3<=2;bcd2<=5;bcd1<=0;bcd0<=9; end
			2510: begin bcd3<=2;bcd2<=5;bcd1<=1;bcd0<=0; end
			2511: begin bcd3<=2;bcd2<=5;bcd1<=1;bcd0<=1; end
			2512: begin bcd3<=2;bcd2<=5;bcd1<=1;bcd0<=2; end
			2513: begin bcd3<=2;bcd2<=5;bcd1<=1;bcd0<=3; end
			2514: begin bcd3<=2;bcd2<=5;bcd1<=1;bcd0<=4; end
			2515: begin bcd3<=2;bcd2<=5;bcd1<=1;bcd0<=5; end
			2516: begin bcd3<=2;bcd2<=5;bcd1<=1;bcd0<=6; end
			2517: begin bcd3<=2;bcd2<=5;bcd1<=1;bcd0<=7; end
			2518: begin bcd3<=2;bcd2<=5;bcd1<=1;bcd0<=8; end
			2519: begin bcd3<=2;bcd2<=5;bcd1<=1;bcd0<=9; end
			2520: begin bcd3<=2;bcd2<=5;bcd1<=2;bcd0<=0; end
			2521: begin bcd3<=2;bcd2<=5;bcd1<=2;bcd0<=1; end
			2522: begin bcd3<=2;bcd2<=5;bcd1<=2;bcd0<=2; end
			2523: begin bcd3<=2;bcd2<=5;bcd1<=2;bcd0<=3; end
			2524: begin bcd3<=2;bcd2<=5;bcd1<=2;bcd0<=4; end
			2525: begin bcd3<=2;bcd2<=5;bcd1<=2;bcd0<=5; end
			2526: begin bcd3<=2;bcd2<=5;bcd1<=2;bcd0<=6; end
			2527: begin bcd3<=2;bcd2<=5;bcd1<=2;bcd0<=7; end
			2528: begin bcd3<=2;bcd2<=5;bcd1<=2;bcd0<=8; end
			2529: begin bcd3<=2;bcd2<=5;bcd1<=2;bcd0<=9; end
			2530: begin bcd3<=2;bcd2<=5;bcd1<=3;bcd0<=0; end
			2531: begin bcd3<=2;bcd2<=5;bcd1<=3;bcd0<=1; end
			2532: begin bcd3<=2;bcd2<=5;bcd1<=3;bcd0<=2; end
			2533: begin bcd3<=2;bcd2<=5;bcd1<=3;bcd0<=3; end
			2534: begin bcd3<=2;bcd2<=5;bcd1<=3;bcd0<=4; end
			2535: begin bcd3<=2;bcd2<=5;bcd1<=3;bcd0<=5; end
			2536: begin bcd3<=2;bcd2<=5;bcd1<=3;bcd0<=6; end
			2537: begin bcd3<=2;bcd2<=5;bcd1<=3;bcd0<=7; end
			2538: begin bcd3<=2;bcd2<=5;bcd1<=3;bcd0<=8; end
			2539: begin bcd3<=2;bcd2<=5;bcd1<=3;bcd0<=9; end
			2540: begin bcd3<=2;bcd2<=5;bcd1<=4;bcd0<=0; end
			2541: begin bcd3<=2;bcd2<=5;bcd1<=4;bcd0<=1; end
			2542: begin bcd3<=2;bcd2<=5;bcd1<=4;bcd0<=2; end
			2543: begin bcd3<=2;bcd2<=5;bcd1<=4;bcd0<=3; end
			2544: begin bcd3<=2;bcd2<=5;bcd1<=4;bcd0<=4; end
			2545: begin bcd3<=2;bcd2<=5;bcd1<=4;bcd0<=5; end
			2546: begin bcd3<=2;bcd2<=5;bcd1<=4;bcd0<=6; end
			2547: begin bcd3<=2;bcd2<=5;bcd1<=4;bcd0<=7; end
			2548: begin bcd3<=2;bcd2<=5;bcd1<=4;bcd0<=8; end
			2549: begin bcd3<=2;bcd2<=5;bcd1<=4;bcd0<=9; end
			2550: begin bcd3<=2;bcd2<=5;bcd1<=5;bcd0<=0; end
			2551: begin bcd3<=2;bcd2<=5;bcd1<=5;bcd0<=1; end
			2552: begin bcd3<=2;bcd2<=5;bcd1<=5;bcd0<=2; end
			2553: begin bcd3<=2;bcd2<=5;bcd1<=5;bcd0<=3; end
			2554: begin bcd3<=2;bcd2<=5;bcd1<=5;bcd0<=4; end
			2555: begin bcd3<=2;bcd2<=5;bcd1<=5;bcd0<=5; end
			2556: begin bcd3<=2;bcd2<=5;bcd1<=5;bcd0<=6; end
			2557: begin bcd3<=2;bcd2<=5;bcd1<=5;bcd0<=7; end
			2558: begin bcd3<=2;bcd2<=5;bcd1<=5;bcd0<=8; end
			2559: begin bcd3<=2;bcd2<=5;bcd1<=5;bcd0<=9; end
			2560: begin bcd3<=2;bcd2<=5;bcd1<=6;bcd0<=0; end
			2561: begin bcd3<=2;bcd2<=5;bcd1<=6;bcd0<=1; end
			2562: begin bcd3<=2;bcd2<=5;bcd1<=6;bcd0<=2; end
			2563: begin bcd3<=2;bcd2<=5;bcd1<=6;bcd0<=3; end
			2564: begin bcd3<=2;bcd2<=5;bcd1<=6;bcd0<=4; end
			2565: begin bcd3<=2;bcd2<=5;bcd1<=6;bcd0<=5; end
			2566: begin bcd3<=2;bcd2<=5;bcd1<=6;bcd0<=6; end
			2567: begin bcd3<=2;bcd2<=5;bcd1<=6;bcd0<=7; end
			2568: begin bcd3<=2;bcd2<=5;bcd1<=6;bcd0<=8; end
			2569: begin bcd3<=2;bcd2<=5;bcd1<=6;bcd0<=9; end
			2570: begin bcd3<=2;bcd2<=5;bcd1<=7;bcd0<=0; end
			2571: begin bcd3<=2;bcd2<=5;bcd1<=7;bcd0<=1; end
			2572: begin bcd3<=2;bcd2<=5;bcd1<=7;bcd0<=2; end
			2573: begin bcd3<=2;bcd2<=5;bcd1<=7;bcd0<=3; end
			2574: begin bcd3<=2;bcd2<=5;bcd1<=7;bcd0<=4; end
			2575: begin bcd3<=2;bcd2<=5;bcd1<=7;bcd0<=5; end
			2576: begin bcd3<=2;bcd2<=5;bcd1<=7;bcd0<=6; end
			2577: begin bcd3<=2;bcd2<=5;bcd1<=7;bcd0<=7; end
			2578: begin bcd3<=2;bcd2<=5;bcd1<=7;bcd0<=8; end
			2579: begin bcd3<=2;bcd2<=5;bcd1<=7;bcd0<=9; end
			2580: begin bcd3<=2;bcd2<=5;bcd1<=8;bcd0<=0; end
			2581: begin bcd3<=2;bcd2<=5;bcd1<=8;bcd0<=1; end
			2582: begin bcd3<=2;bcd2<=5;bcd1<=8;bcd0<=2; end
			2583: begin bcd3<=2;bcd2<=5;bcd1<=8;bcd0<=3; end
			2584: begin bcd3<=2;bcd2<=5;bcd1<=8;bcd0<=4; end
			2585: begin bcd3<=2;bcd2<=5;bcd1<=8;bcd0<=5; end
			2586: begin bcd3<=2;bcd2<=5;bcd1<=8;bcd0<=6; end
			2587: begin bcd3<=2;bcd2<=5;bcd1<=8;bcd0<=7; end
			2588: begin bcd3<=2;bcd2<=5;bcd1<=8;bcd0<=8; end
			2589: begin bcd3<=2;bcd2<=5;bcd1<=8;bcd0<=9; end
			2590: begin bcd3<=2;bcd2<=5;bcd1<=9;bcd0<=0; end
			2591: begin bcd3<=2;bcd2<=5;bcd1<=9;bcd0<=1; end
			2592: begin bcd3<=2;bcd2<=5;bcd1<=9;bcd0<=2; end
			2593: begin bcd3<=2;bcd2<=5;bcd1<=9;bcd0<=3; end
			2594: begin bcd3<=2;bcd2<=5;bcd1<=9;bcd0<=4; end
			2595: begin bcd3<=2;bcd2<=5;bcd1<=9;bcd0<=5; end
			2596: begin bcd3<=2;bcd2<=5;bcd1<=9;bcd0<=6; end
			2597: begin bcd3<=2;bcd2<=5;bcd1<=9;bcd0<=7; end
			2598: begin bcd3<=2;bcd2<=5;bcd1<=9;bcd0<=8; end
			2599: begin bcd3<=2;bcd2<=5;bcd1<=9;bcd0<=9; end
			2600: begin bcd3<=2;bcd2<=6;bcd1<=0;bcd0<=0; end
			2601: begin bcd3<=2;bcd2<=6;bcd1<=0;bcd0<=1; end
			2602: begin bcd3<=2;bcd2<=6;bcd1<=0;bcd0<=2; end
			2603: begin bcd3<=2;bcd2<=6;bcd1<=0;bcd0<=3; end
			2604: begin bcd3<=2;bcd2<=6;bcd1<=0;bcd0<=4; end
			2605: begin bcd3<=2;bcd2<=6;bcd1<=0;bcd0<=5; end
			2606: begin bcd3<=2;bcd2<=6;bcd1<=0;bcd0<=6; end
			2607: begin bcd3<=2;bcd2<=6;bcd1<=0;bcd0<=7; end
			2608: begin bcd3<=2;bcd2<=6;bcd1<=0;bcd0<=8; end
			2609: begin bcd3<=2;bcd2<=6;bcd1<=0;bcd0<=9; end
			2610: begin bcd3<=2;bcd2<=6;bcd1<=1;bcd0<=0; end
			2611: begin bcd3<=2;bcd2<=6;bcd1<=1;bcd0<=1; end
			2612: begin bcd3<=2;bcd2<=6;bcd1<=1;bcd0<=2; end
			2613: begin bcd3<=2;bcd2<=6;bcd1<=1;bcd0<=3; end
			2614: begin bcd3<=2;bcd2<=6;bcd1<=1;bcd0<=4; end
			2615: begin bcd3<=2;bcd2<=6;bcd1<=1;bcd0<=5; end
			2616: begin bcd3<=2;bcd2<=6;bcd1<=1;bcd0<=6; end
			2617: begin bcd3<=2;bcd2<=6;bcd1<=1;bcd0<=7; end
			2618: begin bcd3<=2;bcd2<=6;bcd1<=1;bcd0<=8; end
			2619: begin bcd3<=2;bcd2<=6;bcd1<=1;bcd0<=9; end
			2620: begin bcd3<=2;bcd2<=6;bcd1<=2;bcd0<=0; end
			2621: begin bcd3<=2;bcd2<=6;bcd1<=2;bcd0<=1; end
			2622: begin bcd3<=2;bcd2<=6;bcd1<=2;bcd0<=2; end
			2623: begin bcd3<=2;bcd2<=6;bcd1<=2;bcd0<=3; end
			2624: begin bcd3<=2;bcd2<=6;bcd1<=2;bcd0<=4; end
			2625: begin bcd3<=2;bcd2<=6;bcd1<=2;bcd0<=5; end
			2626: begin bcd3<=2;bcd2<=6;bcd1<=2;bcd0<=6; end
			2627: begin bcd3<=2;bcd2<=6;bcd1<=2;bcd0<=7; end
			2628: begin bcd3<=2;bcd2<=6;bcd1<=2;bcd0<=8; end
			2629: begin bcd3<=2;bcd2<=6;bcd1<=2;bcd0<=9; end
			2630: begin bcd3<=2;bcd2<=6;bcd1<=3;bcd0<=0; end
			2631: begin bcd3<=2;bcd2<=6;bcd1<=3;bcd0<=1; end
			2632: begin bcd3<=2;bcd2<=6;bcd1<=3;bcd0<=2; end
			2633: begin bcd3<=2;bcd2<=6;bcd1<=3;bcd0<=3; end
			2634: begin bcd3<=2;bcd2<=6;bcd1<=3;bcd0<=4; end
			2635: begin bcd3<=2;bcd2<=6;bcd1<=3;bcd0<=5; end
			2636: begin bcd3<=2;bcd2<=6;bcd1<=3;bcd0<=6; end
			2637: begin bcd3<=2;bcd2<=6;bcd1<=3;bcd0<=7; end
			2638: begin bcd3<=2;bcd2<=6;bcd1<=3;bcd0<=8; end
			2639: begin bcd3<=2;bcd2<=6;bcd1<=3;bcd0<=9; end
			2640: begin bcd3<=2;bcd2<=6;bcd1<=4;bcd0<=0; end
			2641: begin bcd3<=2;bcd2<=6;bcd1<=4;bcd0<=1; end
			2642: begin bcd3<=2;bcd2<=6;bcd1<=4;bcd0<=2; end
			2643: begin bcd3<=2;bcd2<=6;bcd1<=4;bcd0<=3; end
			2644: begin bcd3<=2;bcd2<=6;bcd1<=4;bcd0<=4; end
			2645: begin bcd3<=2;bcd2<=6;bcd1<=4;bcd0<=5; end
			2646: begin bcd3<=2;bcd2<=6;bcd1<=4;bcd0<=6; end
			2647: begin bcd3<=2;bcd2<=6;bcd1<=4;bcd0<=7; end
			2648: begin bcd3<=2;bcd2<=6;bcd1<=4;bcd0<=8; end
			2649: begin bcd3<=2;bcd2<=6;bcd1<=4;bcd0<=9; end
			2650: begin bcd3<=2;bcd2<=6;bcd1<=5;bcd0<=0; end
			2651: begin bcd3<=2;bcd2<=6;bcd1<=5;bcd0<=1; end
			2652: begin bcd3<=2;bcd2<=6;bcd1<=5;bcd0<=2; end
			2653: begin bcd3<=2;bcd2<=6;bcd1<=5;bcd0<=3; end
			2654: begin bcd3<=2;bcd2<=6;bcd1<=5;bcd0<=4; end
			2655: begin bcd3<=2;bcd2<=6;bcd1<=5;bcd0<=5; end
			2656: begin bcd3<=2;bcd2<=6;bcd1<=5;bcd0<=6; end
			2657: begin bcd3<=2;bcd2<=6;bcd1<=5;bcd0<=7; end
			2658: begin bcd3<=2;bcd2<=6;bcd1<=5;bcd0<=8; end
			2659: begin bcd3<=2;bcd2<=6;bcd1<=5;bcd0<=9; end
			2660: begin bcd3<=2;bcd2<=6;bcd1<=6;bcd0<=0; end
			2661: begin bcd3<=2;bcd2<=6;bcd1<=6;bcd0<=1; end
			2662: begin bcd3<=2;bcd2<=6;bcd1<=6;bcd0<=2; end
			2663: begin bcd3<=2;bcd2<=6;bcd1<=6;bcd0<=3; end
			2664: begin bcd3<=2;bcd2<=6;bcd1<=6;bcd0<=4; end
			2665: begin bcd3<=2;bcd2<=6;bcd1<=6;bcd0<=5; end
			2666: begin bcd3<=2;bcd2<=6;bcd1<=6;bcd0<=6; end
			2667: begin bcd3<=2;bcd2<=6;bcd1<=6;bcd0<=7; end
			2668: begin bcd3<=2;bcd2<=6;bcd1<=6;bcd0<=8; end
			2669: begin bcd3<=2;bcd2<=6;bcd1<=6;bcd0<=9; end
			2670: begin bcd3<=2;bcd2<=6;bcd1<=7;bcd0<=0; end
			2671: begin bcd3<=2;bcd2<=6;bcd1<=7;bcd0<=1; end
			2672: begin bcd3<=2;bcd2<=6;bcd1<=7;bcd0<=2; end
			2673: begin bcd3<=2;bcd2<=6;bcd1<=7;bcd0<=3; end
			2674: begin bcd3<=2;bcd2<=6;bcd1<=7;bcd0<=4; end
			2675: begin bcd3<=2;bcd2<=6;bcd1<=7;bcd0<=5; end
			2676: begin bcd3<=2;bcd2<=6;bcd1<=7;bcd0<=6; end
			2677: begin bcd3<=2;bcd2<=6;bcd1<=7;bcd0<=7; end
			2678: begin bcd3<=2;bcd2<=6;bcd1<=7;bcd0<=8; end
			2679: begin bcd3<=2;bcd2<=6;bcd1<=7;bcd0<=9; end
			2680: begin bcd3<=2;bcd2<=6;bcd1<=8;bcd0<=0; end
			2681: begin bcd3<=2;bcd2<=6;bcd1<=8;bcd0<=1; end
			2682: begin bcd3<=2;bcd2<=6;bcd1<=8;bcd0<=2; end
			2683: begin bcd3<=2;bcd2<=6;bcd1<=8;bcd0<=3; end
			2684: begin bcd3<=2;bcd2<=6;bcd1<=8;bcd0<=4; end
			2685: begin bcd3<=2;bcd2<=6;bcd1<=8;bcd0<=5; end
			2686: begin bcd3<=2;bcd2<=6;bcd1<=8;bcd0<=6; end
			2687: begin bcd3<=2;bcd2<=6;bcd1<=8;bcd0<=7; end
			2688: begin bcd3<=2;bcd2<=6;bcd1<=8;bcd0<=8; end
			2689: begin bcd3<=2;bcd2<=6;bcd1<=8;bcd0<=9; end
			2690: begin bcd3<=2;bcd2<=6;bcd1<=9;bcd0<=0; end
			2691: begin bcd3<=2;bcd2<=6;bcd1<=9;bcd0<=1; end
			2692: begin bcd3<=2;bcd2<=6;bcd1<=9;bcd0<=2; end
			2693: begin bcd3<=2;bcd2<=6;bcd1<=9;bcd0<=3; end
			2694: begin bcd3<=2;bcd2<=6;bcd1<=9;bcd0<=4; end
			2695: begin bcd3<=2;bcd2<=6;bcd1<=9;bcd0<=5; end
			2696: begin bcd3<=2;bcd2<=6;bcd1<=9;bcd0<=6; end
			2697: begin bcd3<=2;bcd2<=6;bcd1<=9;bcd0<=7; end
			2698: begin bcd3<=2;bcd2<=6;bcd1<=9;bcd0<=8; end
			2699: begin bcd3<=2;bcd2<=6;bcd1<=9;bcd0<=9; end
			2700: begin bcd3<=2;bcd2<=7;bcd1<=0;bcd0<=0; end
			2701: begin bcd3<=2;bcd2<=7;bcd1<=0;bcd0<=1; end
			2702: begin bcd3<=2;bcd2<=7;bcd1<=0;bcd0<=2; end
			2703: begin bcd3<=2;bcd2<=7;bcd1<=0;bcd0<=3; end
			2704: begin bcd3<=2;bcd2<=7;bcd1<=0;bcd0<=4; end
			2705: begin bcd3<=2;bcd2<=7;bcd1<=0;bcd0<=5; end
			2706: begin bcd3<=2;bcd2<=7;bcd1<=0;bcd0<=6; end
			2707: begin bcd3<=2;bcd2<=7;bcd1<=0;bcd0<=7; end
			2708: begin bcd3<=2;bcd2<=7;bcd1<=0;bcd0<=8; end
			2709: begin bcd3<=2;bcd2<=7;bcd1<=0;bcd0<=9; end
			2710: begin bcd3<=2;bcd2<=7;bcd1<=1;bcd0<=0; end
			2711: begin bcd3<=2;bcd2<=7;bcd1<=1;bcd0<=1; end
			2712: begin bcd3<=2;bcd2<=7;bcd1<=1;bcd0<=2; end
			2713: begin bcd3<=2;bcd2<=7;bcd1<=1;bcd0<=3; end
			2714: begin bcd3<=2;bcd2<=7;bcd1<=1;bcd0<=4; end
			2715: begin bcd3<=2;bcd2<=7;bcd1<=1;bcd0<=5; end
			2716: begin bcd3<=2;bcd2<=7;bcd1<=1;bcd0<=6; end
			2717: begin bcd3<=2;bcd2<=7;bcd1<=1;bcd0<=7; end
			2718: begin bcd3<=2;bcd2<=7;bcd1<=1;bcd0<=8; end
			2719: begin bcd3<=2;bcd2<=7;bcd1<=1;bcd0<=9; end
			2720: begin bcd3<=2;bcd2<=7;bcd1<=2;bcd0<=0; end
			2721: begin bcd3<=2;bcd2<=7;bcd1<=2;bcd0<=1; end
			2722: begin bcd3<=2;bcd2<=7;bcd1<=2;bcd0<=2; end
			2723: begin bcd3<=2;bcd2<=7;bcd1<=2;bcd0<=3; end
			2724: begin bcd3<=2;bcd2<=7;bcd1<=2;bcd0<=4; end
			2725: begin bcd3<=2;bcd2<=7;bcd1<=2;bcd0<=5; end
			2726: begin bcd3<=2;bcd2<=7;bcd1<=2;bcd0<=6; end
			2727: begin bcd3<=2;bcd2<=7;bcd1<=2;bcd0<=7; end
			2728: begin bcd3<=2;bcd2<=7;bcd1<=2;bcd0<=8; end
			2729: begin bcd3<=2;bcd2<=7;bcd1<=2;bcd0<=9; end
			2730: begin bcd3<=2;bcd2<=7;bcd1<=3;bcd0<=0; end
			2731: begin bcd3<=2;bcd2<=7;bcd1<=3;bcd0<=1; end
			2732: begin bcd3<=2;bcd2<=7;bcd1<=3;bcd0<=2; end
			2733: begin bcd3<=2;bcd2<=7;bcd1<=3;bcd0<=3; end
			2734: begin bcd3<=2;bcd2<=7;bcd1<=3;bcd0<=4; end
			2735: begin bcd3<=2;bcd2<=7;bcd1<=3;bcd0<=5; end
			2736: begin bcd3<=2;bcd2<=7;bcd1<=3;bcd0<=6; end
			2737: begin bcd3<=2;bcd2<=7;bcd1<=3;bcd0<=7; end
			2738: begin bcd3<=2;bcd2<=7;bcd1<=3;bcd0<=8; end
			2739: begin bcd3<=2;bcd2<=7;bcd1<=3;bcd0<=9; end
			2740: begin bcd3<=2;bcd2<=7;bcd1<=4;bcd0<=0; end
			2741: begin bcd3<=2;bcd2<=7;bcd1<=4;bcd0<=1; end
			2742: begin bcd3<=2;bcd2<=7;bcd1<=4;bcd0<=2; end
			2743: begin bcd3<=2;bcd2<=7;bcd1<=4;bcd0<=3; end
			2744: begin bcd3<=2;bcd2<=7;bcd1<=4;bcd0<=4; end
			2745: begin bcd3<=2;bcd2<=7;bcd1<=4;bcd0<=5; end
			2746: begin bcd3<=2;bcd2<=7;bcd1<=4;bcd0<=6; end
			2747: begin bcd3<=2;bcd2<=7;bcd1<=4;bcd0<=7; end
			2748: begin bcd3<=2;bcd2<=7;bcd1<=4;bcd0<=8; end
			2749: begin bcd3<=2;bcd2<=7;bcd1<=4;bcd0<=9; end
			2750: begin bcd3<=2;bcd2<=7;bcd1<=5;bcd0<=0; end
			2751: begin bcd3<=2;bcd2<=7;bcd1<=5;bcd0<=1; end
			2752: begin bcd3<=2;bcd2<=7;bcd1<=5;bcd0<=2; end
			2753: begin bcd3<=2;bcd2<=7;bcd1<=5;bcd0<=3; end
			2754: begin bcd3<=2;bcd2<=7;bcd1<=5;bcd0<=4; end
			2755: begin bcd3<=2;bcd2<=7;bcd1<=5;bcd0<=5; end
			2756: begin bcd3<=2;bcd2<=7;bcd1<=5;bcd0<=6; end
			2757: begin bcd3<=2;bcd2<=7;bcd1<=5;bcd0<=7; end
			2758: begin bcd3<=2;bcd2<=7;bcd1<=5;bcd0<=8; end
			2759: begin bcd3<=2;bcd2<=7;bcd1<=5;bcd0<=9; end
			2760: begin bcd3<=2;bcd2<=7;bcd1<=6;bcd0<=0; end
			2761: begin bcd3<=2;bcd2<=7;bcd1<=6;bcd0<=1; end
			2762: begin bcd3<=2;bcd2<=7;bcd1<=6;bcd0<=2; end
			2763: begin bcd3<=2;bcd2<=7;bcd1<=6;bcd0<=3; end
			2764: begin bcd3<=2;bcd2<=7;bcd1<=6;bcd0<=4; end
			2765: begin bcd3<=2;bcd2<=7;bcd1<=6;bcd0<=5; end
			2766: begin bcd3<=2;bcd2<=7;bcd1<=6;bcd0<=6; end
			2767: begin bcd3<=2;bcd2<=7;bcd1<=6;bcd0<=7; end
			2768: begin bcd3<=2;bcd2<=7;bcd1<=6;bcd0<=8; end
			2769: begin bcd3<=2;bcd2<=7;bcd1<=6;bcd0<=9; end
			2770: begin bcd3<=2;bcd2<=7;bcd1<=7;bcd0<=0; end
			2771: begin bcd3<=2;bcd2<=7;bcd1<=7;bcd0<=1; end
			2772: begin bcd3<=2;bcd2<=7;bcd1<=7;bcd0<=2; end
			2773: begin bcd3<=2;bcd2<=7;bcd1<=7;bcd0<=3; end
			2774: begin bcd3<=2;bcd2<=7;bcd1<=7;bcd0<=4; end
			2775: begin bcd3<=2;bcd2<=7;bcd1<=7;bcd0<=5; end
			2776: begin bcd3<=2;bcd2<=7;bcd1<=7;bcd0<=6; end
			2777: begin bcd3<=2;bcd2<=7;bcd1<=7;bcd0<=7; end
			2778: begin bcd3<=2;bcd2<=7;bcd1<=7;bcd0<=8; end
			2779: begin bcd3<=2;bcd2<=7;bcd1<=7;bcd0<=9; end
			2780: begin bcd3<=2;bcd2<=7;bcd1<=8;bcd0<=0; end
			2781: begin bcd3<=2;bcd2<=7;bcd1<=8;bcd0<=1; end
			2782: begin bcd3<=2;bcd2<=7;bcd1<=8;bcd0<=2; end
			2783: begin bcd3<=2;bcd2<=7;bcd1<=8;bcd0<=3; end
			2784: begin bcd3<=2;bcd2<=7;bcd1<=8;bcd0<=4; end
			2785: begin bcd3<=2;bcd2<=7;bcd1<=8;bcd0<=5; end
			2786: begin bcd3<=2;bcd2<=7;bcd1<=8;bcd0<=6; end
			2787: begin bcd3<=2;bcd2<=7;bcd1<=8;bcd0<=7; end
			2788: begin bcd3<=2;bcd2<=7;bcd1<=8;bcd0<=8; end
			2789: begin bcd3<=2;bcd2<=7;bcd1<=8;bcd0<=9; end
			2790: begin bcd3<=2;bcd2<=7;bcd1<=9;bcd0<=0; end
			2791: begin bcd3<=2;bcd2<=7;bcd1<=9;bcd0<=1; end
			2792: begin bcd3<=2;bcd2<=7;bcd1<=9;bcd0<=2; end
			2793: begin bcd3<=2;bcd2<=7;bcd1<=9;bcd0<=3; end
			2794: begin bcd3<=2;bcd2<=7;bcd1<=9;bcd0<=4; end
			2795: begin bcd3<=2;bcd2<=7;bcd1<=9;bcd0<=5; end
			2796: begin bcd3<=2;bcd2<=7;bcd1<=9;bcd0<=6; end
			2797: begin bcd3<=2;bcd2<=7;bcd1<=9;bcd0<=7; end
			2798: begin bcd3<=2;bcd2<=7;bcd1<=9;bcd0<=8; end
			2799: begin bcd3<=2;bcd2<=7;bcd1<=9;bcd0<=9; end
			2800: begin bcd3<=2;bcd2<=8;bcd1<=0;bcd0<=0; end
			2801: begin bcd3<=2;bcd2<=8;bcd1<=0;bcd0<=1; end
			2802: begin bcd3<=2;bcd2<=8;bcd1<=0;bcd0<=2; end
			2803: begin bcd3<=2;bcd2<=8;bcd1<=0;bcd0<=3; end
			2804: begin bcd3<=2;bcd2<=8;bcd1<=0;bcd0<=4; end
			2805: begin bcd3<=2;bcd2<=8;bcd1<=0;bcd0<=5; end
			2806: begin bcd3<=2;bcd2<=8;bcd1<=0;bcd0<=6; end
			2807: begin bcd3<=2;bcd2<=8;bcd1<=0;bcd0<=7; end
			2808: begin bcd3<=2;bcd2<=8;bcd1<=0;bcd0<=8; end
			2809: begin bcd3<=2;bcd2<=8;bcd1<=0;bcd0<=9; end
			2810: begin bcd3<=2;bcd2<=8;bcd1<=1;bcd0<=0; end
			2811: begin bcd3<=2;bcd2<=8;bcd1<=1;bcd0<=1; end
			2812: begin bcd3<=2;bcd2<=8;bcd1<=1;bcd0<=2; end
			2813: begin bcd3<=2;bcd2<=8;bcd1<=1;bcd0<=3; end
			2814: begin bcd3<=2;bcd2<=8;bcd1<=1;bcd0<=4; end
			2815: begin bcd3<=2;bcd2<=8;bcd1<=1;bcd0<=5; end
			2816: begin bcd3<=2;bcd2<=8;bcd1<=1;bcd0<=6; end
			2817: begin bcd3<=2;bcd2<=8;bcd1<=1;bcd0<=7; end
			2818: begin bcd3<=2;bcd2<=8;bcd1<=1;bcd0<=8; end
			2819: begin bcd3<=2;bcd2<=8;bcd1<=1;bcd0<=9; end
			2820: begin bcd3<=2;bcd2<=8;bcd1<=2;bcd0<=0; end
			2821: begin bcd3<=2;bcd2<=8;bcd1<=2;bcd0<=1; end
			2822: begin bcd3<=2;bcd2<=8;bcd1<=2;bcd0<=2; end
			2823: begin bcd3<=2;bcd2<=8;bcd1<=2;bcd0<=3; end
			2824: begin bcd3<=2;bcd2<=8;bcd1<=2;bcd0<=4; end
			2825: begin bcd3<=2;bcd2<=8;bcd1<=2;bcd0<=5; end
			2826: begin bcd3<=2;bcd2<=8;bcd1<=2;bcd0<=6; end
			2827: begin bcd3<=2;bcd2<=8;bcd1<=2;bcd0<=7; end
			2828: begin bcd3<=2;bcd2<=8;bcd1<=2;bcd0<=8; end
			2829: begin bcd3<=2;bcd2<=8;bcd1<=2;bcd0<=9; end
			2830: begin bcd3<=2;bcd2<=8;bcd1<=3;bcd0<=0; end
			2831: begin bcd3<=2;bcd2<=8;bcd1<=3;bcd0<=1; end
			2832: begin bcd3<=2;bcd2<=8;bcd1<=3;bcd0<=2; end
			2833: begin bcd3<=2;bcd2<=8;bcd1<=3;bcd0<=3; end
			2834: begin bcd3<=2;bcd2<=8;bcd1<=3;bcd0<=4; end
			2835: begin bcd3<=2;bcd2<=8;bcd1<=3;bcd0<=5; end
			2836: begin bcd3<=2;bcd2<=8;bcd1<=3;bcd0<=6; end
			2837: begin bcd3<=2;bcd2<=8;bcd1<=3;bcd0<=7; end
			2838: begin bcd3<=2;bcd2<=8;bcd1<=3;bcd0<=8; end
			2839: begin bcd3<=2;bcd2<=8;bcd1<=3;bcd0<=9; end
			2840: begin bcd3<=2;bcd2<=8;bcd1<=4;bcd0<=0; end
			2841: begin bcd3<=2;bcd2<=8;bcd1<=4;bcd0<=1; end
			2842: begin bcd3<=2;bcd2<=8;bcd1<=4;bcd0<=2; end
			2843: begin bcd3<=2;bcd2<=8;bcd1<=4;bcd0<=3; end
			2844: begin bcd3<=2;bcd2<=8;bcd1<=4;bcd0<=4; end
			2845: begin bcd3<=2;bcd2<=8;bcd1<=4;bcd0<=5; end
			2846: begin bcd3<=2;bcd2<=8;bcd1<=4;bcd0<=6; end
			2847: begin bcd3<=2;bcd2<=8;bcd1<=4;bcd0<=7; end
			2848: begin bcd3<=2;bcd2<=8;bcd1<=4;bcd0<=8; end
			2849: begin bcd3<=2;bcd2<=8;bcd1<=4;bcd0<=9; end
			2850: begin bcd3<=2;bcd2<=8;bcd1<=5;bcd0<=0; end
			2851: begin bcd3<=2;bcd2<=8;bcd1<=5;bcd0<=1; end
			2852: begin bcd3<=2;bcd2<=8;bcd1<=5;bcd0<=2; end
			2853: begin bcd3<=2;bcd2<=8;bcd1<=5;bcd0<=3; end
			2854: begin bcd3<=2;bcd2<=8;bcd1<=5;bcd0<=4; end
			2855: begin bcd3<=2;bcd2<=8;bcd1<=5;bcd0<=5; end
			2856: begin bcd3<=2;bcd2<=8;bcd1<=5;bcd0<=6; end
			2857: begin bcd3<=2;bcd2<=8;bcd1<=5;bcd0<=7; end
			2858: begin bcd3<=2;bcd2<=8;bcd1<=5;bcd0<=8; end
			2859: begin bcd3<=2;bcd2<=8;bcd1<=5;bcd0<=9; end
			2860: begin bcd3<=2;bcd2<=8;bcd1<=6;bcd0<=0; end
			2861: begin bcd3<=2;bcd2<=8;bcd1<=6;bcd0<=1; end
			2862: begin bcd3<=2;bcd2<=8;bcd1<=6;bcd0<=2; end
			2863: begin bcd3<=2;bcd2<=8;bcd1<=6;bcd0<=3; end
			2864: begin bcd3<=2;bcd2<=8;bcd1<=6;bcd0<=4; end
			2865: begin bcd3<=2;bcd2<=8;bcd1<=6;bcd0<=5; end
			2866: begin bcd3<=2;bcd2<=8;bcd1<=6;bcd0<=6; end
			2867: begin bcd3<=2;bcd2<=8;bcd1<=6;bcd0<=7; end
			2868: begin bcd3<=2;bcd2<=8;bcd1<=6;bcd0<=8; end
			2869: begin bcd3<=2;bcd2<=8;bcd1<=6;bcd0<=9; end
			2870: begin bcd3<=2;bcd2<=8;bcd1<=7;bcd0<=0; end
			2871: begin bcd3<=2;bcd2<=8;bcd1<=7;bcd0<=1; end
			2872: begin bcd3<=2;bcd2<=8;bcd1<=7;bcd0<=2; end
			2873: begin bcd3<=2;bcd2<=8;bcd1<=7;bcd0<=3; end
			2874: begin bcd3<=2;bcd2<=8;bcd1<=7;bcd0<=4; end
			2875: begin bcd3<=2;bcd2<=8;bcd1<=7;bcd0<=5; end
			2876: begin bcd3<=2;bcd2<=8;bcd1<=7;bcd0<=6; end
			2877: begin bcd3<=2;bcd2<=8;bcd1<=7;bcd0<=7; end
			2878: begin bcd3<=2;bcd2<=8;bcd1<=7;bcd0<=8; end
			2879: begin bcd3<=2;bcd2<=8;bcd1<=7;bcd0<=9; end
			2880: begin bcd3<=2;bcd2<=8;bcd1<=8;bcd0<=0; end
			2881: begin bcd3<=2;bcd2<=8;bcd1<=8;bcd0<=1; end
			2882: begin bcd3<=2;bcd2<=8;bcd1<=8;bcd0<=2; end
			2883: begin bcd3<=2;bcd2<=8;bcd1<=8;bcd0<=3; end
			2884: begin bcd3<=2;bcd2<=8;bcd1<=8;bcd0<=4; end
			2885: begin bcd3<=2;bcd2<=8;bcd1<=8;bcd0<=5; end
			2886: begin bcd3<=2;bcd2<=8;bcd1<=8;bcd0<=6; end
			2887: begin bcd3<=2;bcd2<=8;bcd1<=8;bcd0<=7; end
			2888: begin bcd3<=2;bcd2<=8;bcd1<=8;bcd0<=8; end
			2889: begin bcd3<=2;bcd2<=8;bcd1<=8;bcd0<=9; end
			2890: begin bcd3<=2;bcd2<=8;bcd1<=9;bcd0<=0; end
			2891: begin bcd3<=2;bcd2<=8;bcd1<=9;bcd0<=1; end
			2892: begin bcd3<=2;bcd2<=8;bcd1<=9;bcd0<=2; end
			2893: begin bcd3<=2;bcd2<=8;bcd1<=9;bcd0<=3; end
			2894: begin bcd3<=2;bcd2<=8;bcd1<=9;bcd0<=4; end
			2895: begin bcd3<=2;bcd2<=8;bcd1<=9;bcd0<=5; end
			2896: begin bcd3<=2;bcd2<=8;bcd1<=9;bcd0<=6; end
			2897: begin bcd3<=2;bcd2<=8;bcd1<=9;bcd0<=7; end
			2898: begin bcd3<=2;bcd2<=8;bcd1<=9;bcd0<=8; end
			2899: begin bcd3<=2;bcd2<=8;bcd1<=9;bcd0<=9; end
			2900: begin bcd3<=2;bcd2<=9;bcd1<=0;bcd0<=0; end
			2901: begin bcd3<=2;bcd2<=9;bcd1<=0;bcd0<=1; end
			2902: begin bcd3<=2;bcd2<=9;bcd1<=0;bcd0<=2; end
			2903: begin bcd3<=2;bcd2<=9;bcd1<=0;bcd0<=3; end
			2904: begin bcd3<=2;bcd2<=9;bcd1<=0;bcd0<=4; end
			2905: begin bcd3<=2;bcd2<=9;bcd1<=0;bcd0<=5; end
			2906: begin bcd3<=2;bcd2<=9;bcd1<=0;bcd0<=6; end
			2907: begin bcd3<=2;bcd2<=9;bcd1<=0;bcd0<=7; end
			2908: begin bcd3<=2;bcd2<=9;bcd1<=0;bcd0<=8; end
			2909: begin bcd3<=2;bcd2<=9;bcd1<=0;bcd0<=9; end
			2910: begin bcd3<=2;bcd2<=9;bcd1<=1;bcd0<=0; end
			2911: begin bcd3<=2;bcd2<=9;bcd1<=1;bcd0<=1; end
			2912: begin bcd3<=2;bcd2<=9;bcd1<=1;bcd0<=2; end
			2913: begin bcd3<=2;bcd2<=9;bcd1<=1;bcd0<=3; end
			2914: begin bcd3<=2;bcd2<=9;bcd1<=1;bcd0<=4; end
			2915: begin bcd3<=2;bcd2<=9;bcd1<=1;bcd0<=5; end
			2916: begin bcd3<=2;bcd2<=9;bcd1<=1;bcd0<=6; end
			2917: begin bcd3<=2;bcd2<=9;bcd1<=1;bcd0<=7; end
			2918: begin bcd3<=2;bcd2<=9;bcd1<=1;bcd0<=8; end
			2919: begin bcd3<=2;bcd2<=9;bcd1<=1;bcd0<=9; end
			2920: begin bcd3<=2;bcd2<=9;bcd1<=2;bcd0<=0; end
			2921: begin bcd3<=2;bcd2<=9;bcd1<=2;bcd0<=1; end
			2922: begin bcd3<=2;bcd2<=9;bcd1<=2;bcd0<=2; end
			2923: begin bcd3<=2;bcd2<=9;bcd1<=2;bcd0<=3; end
			2924: begin bcd3<=2;bcd2<=9;bcd1<=2;bcd0<=4; end
			2925: begin bcd3<=2;bcd2<=9;bcd1<=2;bcd0<=5; end
			2926: begin bcd3<=2;bcd2<=9;bcd1<=2;bcd0<=6; end
			2927: begin bcd3<=2;bcd2<=9;bcd1<=2;bcd0<=7; end
			2928: begin bcd3<=2;bcd2<=9;bcd1<=2;bcd0<=8; end
			2929: begin bcd3<=2;bcd2<=9;bcd1<=2;bcd0<=9; end
			2930: begin bcd3<=2;bcd2<=9;bcd1<=3;bcd0<=0; end
			2931: begin bcd3<=2;bcd2<=9;bcd1<=3;bcd0<=1; end
			2932: begin bcd3<=2;bcd2<=9;bcd1<=3;bcd0<=2; end
			2933: begin bcd3<=2;bcd2<=9;bcd1<=3;bcd0<=3; end
			2934: begin bcd3<=2;bcd2<=9;bcd1<=3;bcd0<=4; end
			2935: begin bcd3<=2;bcd2<=9;bcd1<=3;bcd0<=5; end
			2936: begin bcd3<=2;bcd2<=9;bcd1<=3;bcd0<=6; end
			2937: begin bcd3<=2;bcd2<=9;bcd1<=3;bcd0<=7; end
			2938: begin bcd3<=2;bcd2<=9;bcd1<=3;bcd0<=8; end
			2939: begin bcd3<=2;bcd2<=9;bcd1<=3;bcd0<=9; end
			2940: begin bcd3<=2;bcd2<=9;bcd1<=4;bcd0<=0; end
			2941: begin bcd3<=2;bcd2<=9;bcd1<=4;bcd0<=1; end
			2942: begin bcd3<=2;bcd2<=9;bcd1<=4;bcd0<=2; end
			2943: begin bcd3<=2;bcd2<=9;bcd1<=4;bcd0<=3; end
			2944: begin bcd3<=2;bcd2<=9;bcd1<=4;bcd0<=4; end
			2945: begin bcd3<=2;bcd2<=9;bcd1<=4;bcd0<=5; end
			2946: begin bcd3<=2;bcd2<=9;bcd1<=4;bcd0<=6; end
			2947: begin bcd3<=2;bcd2<=9;bcd1<=4;bcd0<=7; end
			2948: begin bcd3<=2;bcd2<=9;bcd1<=4;bcd0<=8; end
			2949: begin bcd3<=2;bcd2<=9;bcd1<=4;bcd0<=9; end
			2950: begin bcd3<=2;bcd2<=9;bcd1<=5;bcd0<=0; end
			2951: begin bcd3<=2;bcd2<=9;bcd1<=5;bcd0<=1; end
			2952: begin bcd3<=2;bcd2<=9;bcd1<=5;bcd0<=2; end
			2953: begin bcd3<=2;bcd2<=9;bcd1<=5;bcd0<=3; end
			2954: begin bcd3<=2;bcd2<=9;bcd1<=5;bcd0<=4; end
			2955: begin bcd3<=2;bcd2<=9;bcd1<=5;bcd0<=5; end
			2956: begin bcd3<=2;bcd2<=9;bcd1<=5;bcd0<=6; end
			2957: begin bcd3<=2;bcd2<=9;bcd1<=5;bcd0<=7; end
			2958: begin bcd3<=2;bcd2<=9;bcd1<=5;bcd0<=8; end
			2959: begin bcd3<=2;bcd2<=9;bcd1<=5;bcd0<=9; end
			2960: begin bcd3<=2;bcd2<=9;bcd1<=6;bcd0<=0; end
			2961: begin bcd3<=2;bcd2<=9;bcd1<=6;bcd0<=1; end
			2962: begin bcd3<=2;bcd2<=9;bcd1<=6;bcd0<=2; end
			2963: begin bcd3<=2;bcd2<=9;bcd1<=6;bcd0<=3; end
			2964: begin bcd3<=2;bcd2<=9;bcd1<=6;bcd0<=4; end
			2965: begin bcd3<=2;bcd2<=9;bcd1<=6;bcd0<=5; end
			2966: begin bcd3<=2;bcd2<=9;bcd1<=6;bcd0<=6; end
			2967: begin bcd3<=2;bcd2<=9;bcd1<=6;bcd0<=7; end
			2968: begin bcd3<=2;bcd2<=9;bcd1<=6;bcd0<=8; end
			2969: begin bcd3<=2;bcd2<=9;bcd1<=6;bcd0<=9; end
			2970: begin bcd3<=2;bcd2<=9;bcd1<=7;bcd0<=0; end
			2971: begin bcd3<=2;bcd2<=9;bcd1<=7;bcd0<=1; end
			2972: begin bcd3<=2;bcd2<=9;bcd1<=7;bcd0<=2; end
			2973: begin bcd3<=2;bcd2<=9;bcd1<=7;bcd0<=3; end
			2974: begin bcd3<=2;bcd2<=9;bcd1<=7;bcd0<=4; end
			2975: begin bcd3<=2;bcd2<=9;bcd1<=7;bcd0<=5; end
			2976: begin bcd3<=2;bcd2<=9;bcd1<=7;bcd0<=6; end
			2977: begin bcd3<=2;bcd2<=9;bcd1<=7;bcd0<=7; end
			2978: begin bcd3<=2;bcd2<=9;bcd1<=7;bcd0<=8; end
			2979: begin bcd3<=2;bcd2<=9;bcd1<=7;bcd0<=9; end
			2980: begin bcd3<=2;bcd2<=9;bcd1<=8;bcd0<=0; end
			2981: begin bcd3<=2;bcd2<=9;bcd1<=8;bcd0<=1; end
			2982: begin bcd3<=2;bcd2<=9;bcd1<=8;bcd0<=2; end
			2983: begin bcd3<=2;bcd2<=9;bcd1<=8;bcd0<=3; end
			2984: begin bcd3<=2;bcd2<=9;bcd1<=8;bcd0<=4; end
			2985: begin bcd3<=2;bcd2<=9;bcd1<=8;bcd0<=5; end
			2986: begin bcd3<=2;bcd2<=9;bcd1<=8;bcd0<=6; end
			2987: begin bcd3<=2;bcd2<=9;bcd1<=8;bcd0<=7; end
			2988: begin bcd3<=2;bcd2<=9;bcd1<=8;bcd0<=8; end
			2989: begin bcd3<=2;bcd2<=9;bcd1<=8;bcd0<=9; end
			2990: begin bcd3<=2;bcd2<=9;bcd1<=9;bcd0<=0; end
			2991: begin bcd3<=2;bcd2<=9;bcd1<=9;bcd0<=1; end
			2992: begin bcd3<=2;bcd2<=9;bcd1<=9;bcd0<=2; end
			2993: begin bcd3<=2;bcd2<=9;bcd1<=9;bcd0<=3; end
			2994: begin bcd3<=2;bcd2<=9;bcd1<=9;bcd0<=4; end
			2995: begin bcd3<=2;bcd2<=9;bcd1<=9;bcd0<=5; end
			2996: begin bcd3<=2;bcd2<=9;bcd1<=9;bcd0<=6; end
			2997: begin bcd3<=2;bcd2<=9;bcd1<=9;bcd0<=7; end
			2998: begin bcd3<=2;bcd2<=9;bcd1<=9;bcd0<=8; end
			2999: begin bcd3<=2;bcd2<=9;bcd1<=9;bcd0<=9; end
			3000: begin bcd3<=3;bcd2<=0;bcd1<=0;bcd0<=0; end
			3001: begin bcd3<=3;bcd2<=0;bcd1<=0;bcd0<=1; end
			3002: begin bcd3<=3;bcd2<=0;bcd1<=0;bcd0<=2; end
			3003: begin bcd3<=3;bcd2<=0;bcd1<=0;bcd0<=3; end
			3004: begin bcd3<=3;bcd2<=0;bcd1<=0;bcd0<=4; end
			3005: begin bcd3<=3;bcd2<=0;bcd1<=0;bcd0<=5; end
			3006: begin bcd3<=3;bcd2<=0;bcd1<=0;bcd0<=6; end
			3007: begin bcd3<=3;bcd2<=0;bcd1<=0;bcd0<=7; end
			3008: begin bcd3<=3;bcd2<=0;bcd1<=0;bcd0<=8; end
			3009: begin bcd3<=3;bcd2<=0;bcd1<=0;bcd0<=9; end
			3010: begin bcd3<=3;bcd2<=0;bcd1<=1;bcd0<=0; end
			3011: begin bcd3<=3;bcd2<=0;bcd1<=1;bcd0<=1; end
			3012: begin bcd3<=3;bcd2<=0;bcd1<=1;bcd0<=2; end
			3013: begin bcd3<=3;bcd2<=0;bcd1<=1;bcd0<=3; end
			3014: begin bcd3<=3;bcd2<=0;bcd1<=1;bcd0<=4; end
			3015: begin bcd3<=3;bcd2<=0;bcd1<=1;bcd0<=5; end
			3016: begin bcd3<=3;bcd2<=0;bcd1<=1;bcd0<=6; end
			3017: begin bcd3<=3;bcd2<=0;bcd1<=1;bcd0<=7; end
			3018: begin bcd3<=3;bcd2<=0;bcd1<=1;bcd0<=8; end
			3019: begin bcd3<=3;bcd2<=0;bcd1<=1;bcd0<=9; end
			3020: begin bcd3<=3;bcd2<=0;bcd1<=2;bcd0<=0; end
			3021: begin bcd3<=3;bcd2<=0;bcd1<=2;bcd0<=1; end
			3022: begin bcd3<=3;bcd2<=0;bcd1<=2;bcd0<=2; end
			3023: begin bcd3<=3;bcd2<=0;bcd1<=2;bcd0<=3; end
			3024: begin bcd3<=3;bcd2<=0;bcd1<=2;bcd0<=4; end
			3025: begin bcd3<=3;bcd2<=0;bcd1<=2;bcd0<=5; end
			3026: begin bcd3<=3;bcd2<=0;bcd1<=2;bcd0<=6; end
			3027: begin bcd3<=3;bcd2<=0;bcd1<=2;bcd0<=7; end
			3028: begin bcd3<=3;bcd2<=0;bcd1<=2;bcd0<=8; end
			3029: begin bcd3<=3;bcd2<=0;bcd1<=2;bcd0<=9; end
			3030: begin bcd3<=3;bcd2<=0;bcd1<=3;bcd0<=0; end
			3031: begin bcd3<=3;bcd2<=0;bcd1<=3;bcd0<=1; end
			3032: begin bcd3<=3;bcd2<=0;bcd1<=3;bcd0<=2; end
			3033: begin bcd3<=3;bcd2<=0;bcd1<=3;bcd0<=3; end
			3034: begin bcd3<=3;bcd2<=0;bcd1<=3;bcd0<=4; end
			3035: begin bcd3<=3;bcd2<=0;bcd1<=3;bcd0<=5; end
			3036: begin bcd3<=3;bcd2<=0;bcd1<=3;bcd0<=6; end
			3037: begin bcd3<=3;bcd2<=0;bcd1<=3;bcd0<=7; end
			3038: begin bcd3<=3;bcd2<=0;bcd1<=3;bcd0<=8; end
			3039: begin bcd3<=3;bcd2<=0;bcd1<=3;bcd0<=9; end
			3040: begin bcd3<=3;bcd2<=0;bcd1<=4;bcd0<=0; end
			3041: begin bcd3<=3;bcd2<=0;bcd1<=4;bcd0<=1; end
			3042: begin bcd3<=3;bcd2<=0;bcd1<=4;bcd0<=2; end
			3043: begin bcd3<=3;bcd2<=0;bcd1<=4;bcd0<=3; end
			3044: begin bcd3<=3;bcd2<=0;bcd1<=4;bcd0<=4; end
			3045: begin bcd3<=3;bcd2<=0;bcd1<=4;bcd0<=5; end
			3046: begin bcd3<=3;bcd2<=0;bcd1<=4;bcd0<=6; end
			3047: begin bcd3<=3;bcd2<=0;bcd1<=4;bcd0<=7; end
			3048: begin bcd3<=3;bcd2<=0;bcd1<=4;bcd0<=8; end
			3049: begin bcd3<=3;bcd2<=0;bcd1<=4;bcd0<=9; end
			3050: begin bcd3<=3;bcd2<=0;bcd1<=5;bcd0<=0; end
			3051: begin bcd3<=3;bcd2<=0;bcd1<=5;bcd0<=1; end
			3052: begin bcd3<=3;bcd2<=0;bcd1<=5;bcd0<=2; end
			3053: begin bcd3<=3;bcd2<=0;bcd1<=5;bcd0<=3; end
			3054: begin bcd3<=3;bcd2<=0;bcd1<=5;bcd0<=4; end
			3055: begin bcd3<=3;bcd2<=0;bcd1<=5;bcd0<=5; end
			3056: begin bcd3<=3;bcd2<=0;bcd1<=5;bcd0<=6; end
			3057: begin bcd3<=3;bcd2<=0;bcd1<=5;bcd0<=7; end
			3058: begin bcd3<=3;bcd2<=0;bcd1<=5;bcd0<=8; end
			3059: begin bcd3<=3;bcd2<=0;bcd1<=5;bcd0<=9; end
			3060: begin bcd3<=3;bcd2<=0;bcd1<=6;bcd0<=0; end
			3061: begin bcd3<=3;bcd2<=0;bcd1<=6;bcd0<=1; end
			3062: begin bcd3<=3;bcd2<=0;bcd1<=6;bcd0<=2; end
			3063: begin bcd3<=3;bcd2<=0;bcd1<=6;bcd0<=3; end
			3064: begin bcd3<=3;bcd2<=0;bcd1<=6;bcd0<=4; end
			3065: begin bcd3<=3;bcd2<=0;bcd1<=6;bcd0<=5; end
			3066: begin bcd3<=3;bcd2<=0;bcd1<=6;bcd0<=6; end
			3067: begin bcd3<=3;bcd2<=0;bcd1<=6;bcd0<=7; end
			3068: begin bcd3<=3;bcd2<=0;bcd1<=6;bcd0<=8; end
			3069: begin bcd3<=3;bcd2<=0;bcd1<=6;bcd0<=9; end
			3070: begin bcd3<=3;bcd2<=0;bcd1<=7;bcd0<=0; end
			3071: begin bcd3<=3;bcd2<=0;bcd1<=7;bcd0<=1; end
			3072: begin bcd3<=3;bcd2<=0;bcd1<=7;bcd0<=2; end
			3073: begin bcd3<=3;bcd2<=0;bcd1<=7;bcd0<=3; end
			3074: begin bcd3<=3;bcd2<=0;bcd1<=7;bcd0<=4; end
			3075: begin bcd3<=3;bcd2<=0;bcd1<=7;bcd0<=5; end
			3076: begin bcd3<=3;bcd2<=0;bcd1<=7;bcd0<=6; end
			3077: begin bcd3<=3;bcd2<=0;bcd1<=7;bcd0<=7; end
			3078: begin bcd3<=3;bcd2<=0;bcd1<=7;bcd0<=8; end
			3079: begin bcd3<=3;bcd2<=0;bcd1<=7;bcd0<=9; end
			3080: begin bcd3<=3;bcd2<=0;bcd1<=8;bcd0<=0; end
			3081: begin bcd3<=3;bcd2<=0;bcd1<=8;bcd0<=1; end
			3082: begin bcd3<=3;bcd2<=0;bcd1<=8;bcd0<=2; end
			3083: begin bcd3<=3;bcd2<=0;bcd1<=8;bcd0<=3; end
			3084: begin bcd3<=3;bcd2<=0;bcd1<=8;bcd0<=4; end
			3085: begin bcd3<=3;bcd2<=0;bcd1<=8;bcd0<=5; end
			3086: begin bcd3<=3;bcd2<=0;bcd1<=8;bcd0<=6; end
			3087: begin bcd3<=3;bcd2<=0;bcd1<=8;bcd0<=7; end
			3088: begin bcd3<=3;bcd2<=0;bcd1<=8;bcd0<=8; end
			3089: begin bcd3<=3;bcd2<=0;bcd1<=8;bcd0<=9; end
			3090: begin bcd3<=3;bcd2<=0;bcd1<=9;bcd0<=0; end
			3091: begin bcd3<=3;bcd2<=0;bcd1<=9;bcd0<=1; end
			3092: begin bcd3<=3;bcd2<=0;bcd1<=9;bcd0<=2; end
			3093: begin bcd3<=3;bcd2<=0;bcd1<=9;bcd0<=3; end
			3094: begin bcd3<=3;bcd2<=0;bcd1<=9;bcd0<=4; end
			3095: begin bcd3<=3;bcd2<=0;bcd1<=9;bcd0<=5; end
			3096: begin bcd3<=3;bcd2<=0;bcd1<=9;bcd0<=6; end
			3097: begin bcd3<=3;bcd2<=0;bcd1<=9;bcd0<=7; end
			3098: begin bcd3<=3;bcd2<=0;bcd1<=9;bcd0<=8; end
			3099: begin bcd3<=3;bcd2<=0;bcd1<=9;bcd0<=9; end
			3100: begin bcd3<=3;bcd2<=1;bcd1<=0;bcd0<=0; end
			3101: begin bcd3<=3;bcd2<=1;bcd1<=0;bcd0<=1; end
			3102: begin bcd3<=3;bcd2<=1;bcd1<=0;bcd0<=2; end
			3103: begin bcd3<=3;bcd2<=1;bcd1<=0;bcd0<=3; end
			3104: begin bcd3<=3;bcd2<=1;bcd1<=0;bcd0<=4; end
			3105: begin bcd3<=3;bcd2<=1;bcd1<=0;bcd0<=5; end
			3106: begin bcd3<=3;bcd2<=1;bcd1<=0;bcd0<=6; end
			3107: begin bcd3<=3;bcd2<=1;bcd1<=0;bcd0<=7; end
			3108: begin bcd3<=3;bcd2<=1;bcd1<=0;bcd0<=8; end
			3109: begin bcd3<=3;bcd2<=1;bcd1<=0;bcd0<=9; end
			3110: begin bcd3<=3;bcd2<=1;bcd1<=1;bcd0<=0; end
			3111: begin bcd3<=3;bcd2<=1;bcd1<=1;bcd0<=1; end
			3112: begin bcd3<=3;bcd2<=1;bcd1<=1;bcd0<=2; end
			3113: begin bcd3<=3;bcd2<=1;bcd1<=1;bcd0<=3; end
			3114: begin bcd3<=3;bcd2<=1;bcd1<=1;bcd0<=4; end
			3115: begin bcd3<=3;bcd2<=1;bcd1<=1;bcd0<=5; end
			3116: begin bcd3<=3;bcd2<=1;bcd1<=1;bcd0<=6; end
			3117: begin bcd3<=3;bcd2<=1;bcd1<=1;bcd0<=7; end
			3118: begin bcd3<=3;bcd2<=1;bcd1<=1;bcd0<=8; end
			3119: begin bcd3<=3;bcd2<=1;bcd1<=1;bcd0<=9; end
			3120: begin bcd3<=3;bcd2<=1;bcd1<=2;bcd0<=0; end
			3121: begin bcd3<=3;bcd2<=1;bcd1<=2;bcd0<=1; end
			3122: begin bcd3<=3;bcd2<=1;bcd1<=2;bcd0<=2; end
			3123: begin bcd3<=3;bcd2<=1;bcd1<=2;bcd0<=3; end
			3124: begin bcd3<=3;bcd2<=1;bcd1<=2;bcd0<=4; end
			3125: begin bcd3<=3;bcd2<=1;bcd1<=2;bcd0<=5; end
			3126: begin bcd3<=3;bcd2<=1;bcd1<=2;bcd0<=6; end
			3127: begin bcd3<=3;bcd2<=1;bcd1<=2;bcd0<=7; end
			3128: begin bcd3<=3;bcd2<=1;bcd1<=2;bcd0<=8; end
			3129: begin bcd3<=3;bcd2<=1;bcd1<=2;bcd0<=9; end
			3130: begin bcd3<=3;bcd2<=1;bcd1<=3;bcd0<=0; end
			3131: begin bcd3<=3;bcd2<=1;bcd1<=3;bcd0<=1; end
			3132: begin bcd3<=3;bcd2<=1;bcd1<=3;bcd0<=2; end
			3133: begin bcd3<=3;bcd2<=1;bcd1<=3;bcd0<=3; end
			3134: begin bcd3<=3;bcd2<=1;bcd1<=3;bcd0<=4; end
			3135: begin bcd3<=3;bcd2<=1;bcd1<=3;bcd0<=5; end
			3136: begin bcd3<=3;bcd2<=1;bcd1<=3;bcd0<=6; end
			3137: begin bcd3<=3;bcd2<=1;bcd1<=3;bcd0<=7; end
			3138: begin bcd3<=3;bcd2<=1;bcd1<=3;bcd0<=8; end
			3139: begin bcd3<=3;bcd2<=1;bcd1<=3;bcd0<=9; end
			3140: begin bcd3<=3;bcd2<=1;bcd1<=4;bcd0<=0; end
			3141: begin bcd3<=3;bcd2<=1;bcd1<=4;bcd0<=1; end
			3142: begin bcd3<=3;bcd2<=1;bcd1<=4;bcd0<=2; end
			3143: begin bcd3<=3;bcd2<=1;bcd1<=4;bcd0<=3; end
			3144: begin bcd3<=3;bcd2<=1;bcd1<=4;bcd0<=4; end
			3145: begin bcd3<=3;bcd2<=1;bcd1<=4;bcd0<=5; end
			3146: begin bcd3<=3;bcd2<=1;bcd1<=4;bcd0<=6; end
			3147: begin bcd3<=3;bcd2<=1;bcd1<=4;bcd0<=7; end
			3148: begin bcd3<=3;bcd2<=1;bcd1<=4;bcd0<=8; end
			3149: begin bcd3<=3;bcd2<=1;bcd1<=4;bcd0<=9; end
			3150: begin bcd3<=3;bcd2<=1;bcd1<=5;bcd0<=0; end
			3151: begin bcd3<=3;bcd2<=1;bcd1<=5;bcd0<=1; end
			3152: begin bcd3<=3;bcd2<=1;bcd1<=5;bcd0<=2; end
			3153: begin bcd3<=3;bcd2<=1;bcd1<=5;bcd0<=3; end
			3154: begin bcd3<=3;bcd2<=1;bcd1<=5;bcd0<=4; end
			3155: begin bcd3<=3;bcd2<=1;bcd1<=5;bcd0<=5; end
			3156: begin bcd3<=3;bcd2<=1;bcd1<=5;bcd0<=6; end
			3157: begin bcd3<=3;bcd2<=1;bcd1<=5;bcd0<=7; end
			3158: begin bcd3<=3;bcd2<=1;bcd1<=5;bcd0<=8; end
			3159: begin bcd3<=3;bcd2<=1;bcd1<=5;bcd0<=9; end
			3160: begin bcd3<=3;bcd2<=1;bcd1<=6;bcd0<=0; end
			3161: begin bcd3<=3;bcd2<=1;bcd1<=6;bcd0<=1; end
			3162: begin bcd3<=3;bcd2<=1;bcd1<=6;bcd0<=2; end
			3163: begin bcd3<=3;bcd2<=1;bcd1<=6;bcd0<=3; end
			3164: begin bcd3<=3;bcd2<=1;bcd1<=6;bcd0<=4; end
			3165: begin bcd3<=3;bcd2<=1;bcd1<=6;bcd0<=5; end
			3166: begin bcd3<=3;bcd2<=1;bcd1<=6;bcd0<=6; end
			3167: begin bcd3<=3;bcd2<=1;bcd1<=6;bcd0<=7; end
			3168: begin bcd3<=3;bcd2<=1;bcd1<=6;bcd0<=8; end
			3169: begin bcd3<=3;bcd2<=1;bcd1<=6;bcd0<=9; end
			3170: begin bcd3<=3;bcd2<=1;bcd1<=7;bcd0<=0; end
			3171: begin bcd3<=3;bcd2<=1;bcd1<=7;bcd0<=1; end
			3172: begin bcd3<=3;bcd2<=1;bcd1<=7;bcd0<=2; end
			3173: begin bcd3<=3;bcd2<=1;bcd1<=7;bcd0<=3; end
			3174: begin bcd3<=3;bcd2<=1;bcd1<=7;bcd0<=4; end
			3175: begin bcd3<=3;bcd2<=1;bcd1<=7;bcd0<=5; end
			3176: begin bcd3<=3;bcd2<=1;bcd1<=7;bcd0<=6; end
			3177: begin bcd3<=3;bcd2<=1;bcd1<=7;bcd0<=7; end
			3178: begin bcd3<=3;bcd2<=1;bcd1<=7;bcd0<=8; end
			3179: begin bcd3<=3;bcd2<=1;bcd1<=7;bcd0<=9; end
			3180: begin bcd3<=3;bcd2<=1;bcd1<=8;bcd0<=0; end
			3181: begin bcd3<=3;bcd2<=1;bcd1<=8;bcd0<=1; end
			3182: begin bcd3<=3;bcd2<=1;bcd1<=8;bcd0<=2; end
			3183: begin bcd3<=3;bcd2<=1;bcd1<=8;bcd0<=3; end
			3184: begin bcd3<=3;bcd2<=1;bcd1<=8;bcd0<=4; end
			3185: begin bcd3<=3;bcd2<=1;bcd1<=8;bcd0<=5; end
			3186: begin bcd3<=3;bcd2<=1;bcd1<=8;bcd0<=6; end
			3187: begin bcd3<=3;bcd2<=1;bcd1<=8;bcd0<=7; end
			3188: begin bcd3<=3;bcd2<=1;bcd1<=8;bcd0<=8; end
			3189: begin bcd3<=3;bcd2<=1;bcd1<=8;bcd0<=9; end
			3190: begin bcd3<=3;bcd2<=1;bcd1<=9;bcd0<=0; end
			3191: begin bcd3<=3;bcd2<=1;bcd1<=9;bcd0<=1; end
			3192: begin bcd3<=3;bcd2<=1;bcd1<=9;bcd0<=2; end
			3193: begin bcd3<=3;bcd2<=1;bcd1<=9;bcd0<=3; end
			3194: begin bcd3<=3;bcd2<=1;bcd1<=9;bcd0<=4; end
			3195: begin bcd3<=3;bcd2<=1;bcd1<=9;bcd0<=5; end
			3196: begin bcd3<=3;bcd2<=1;bcd1<=9;bcd0<=6; end
			3197: begin bcd3<=3;bcd2<=1;bcd1<=9;bcd0<=7; end
			3198: begin bcd3<=3;bcd2<=1;bcd1<=9;bcd0<=8; end
			3199: begin bcd3<=3;bcd2<=1;bcd1<=9;bcd0<=9; end
			3200: begin bcd3<=3;bcd2<=2;bcd1<=0;bcd0<=0; end
			3201: begin bcd3<=3;bcd2<=2;bcd1<=0;bcd0<=1; end
			3202: begin bcd3<=3;bcd2<=2;bcd1<=0;bcd0<=2; end
			3203: begin bcd3<=3;bcd2<=2;bcd1<=0;bcd0<=3; end
			3204: begin bcd3<=3;bcd2<=2;bcd1<=0;bcd0<=4; end
			3205: begin bcd3<=3;bcd2<=2;bcd1<=0;bcd0<=5; end
			3206: begin bcd3<=3;bcd2<=2;bcd1<=0;bcd0<=6; end
			3207: begin bcd3<=3;bcd2<=2;bcd1<=0;bcd0<=7; end
			3208: begin bcd3<=3;bcd2<=2;bcd1<=0;bcd0<=8; end
			3209: begin bcd3<=3;bcd2<=2;bcd1<=0;bcd0<=9; end
			3210: begin bcd3<=3;bcd2<=2;bcd1<=1;bcd0<=0; end
			3211: begin bcd3<=3;bcd2<=2;bcd1<=1;bcd0<=1; end
			3212: begin bcd3<=3;bcd2<=2;bcd1<=1;bcd0<=2; end
			3213: begin bcd3<=3;bcd2<=2;bcd1<=1;bcd0<=3; end
			3214: begin bcd3<=3;bcd2<=2;bcd1<=1;bcd0<=4; end
			3215: begin bcd3<=3;bcd2<=2;bcd1<=1;bcd0<=5; end
			3216: begin bcd3<=3;bcd2<=2;bcd1<=1;bcd0<=6; end
			3217: begin bcd3<=3;bcd2<=2;bcd1<=1;bcd0<=7; end
			3218: begin bcd3<=3;bcd2<=2;bcd1<=1;bcd0<=8; end
			3219: begin bcd3<=3;bcd2<=2;bcd1<=1;bcd0<=9; end
			3220: begin bcd3<=3;bcd2<=2;bcd1<=2;bcd0<=0; end
			3221: begin bcd3<=3;bcd2<=2;bcd1<=2;bcd0<=1; end
			3222: begin bcd3<=3;bcd2<=2;bcd1<=2;bcd0<=2; end
			3223: begin bcd3<=3;bcd2<=2;bcd1<=2;bcd0<=3; end
			3224: begin bcd3<=3;bcd2<=2;bcd1<=2;bcd0<=4; end
			3225: begin bcd3<=3;bcd2<=2;bcd1<=2;bcd0<=5; end
			3226: begin bcd3<=3;bcd2<=2;bcd1<=2;bcd0<=6; end
			3227: begin bcd3<=3;bcd2<=2;bcd1<=2;bcd0<=7; end
			3228: begin bcd3<=3;bcd2<=2;bcd1<=2;bcd0<=8; end
			3229: begin bcd3<=3;bcd2<=2;bcd1<=2;bcd0<=9; end
			3230: begin bcd3<=3;bcd2<=2;bcd1<=3;bcd0<=0; end
			3231: begin bcd3<=3;bcd2<=2;bcd1<=3;bcd0<=1; end
			3232: begin bcd3<=3;bcd2<=2;bcd1<=3;bcd0<=2; end
			3233: begin bcd3<=3;bcd2<=2;bcd1<=3;bcd0<=3; end
			3234: begin bcd3<=3;bcd2<=2;bcd1<=3;bcd0<=4; end
			3235: begin bcd3<=3;bcd2<=2;bcd1<=3;bcd0<=5; end
			3236: begin bcd3<=3;bcd2<=2;bcd1<=3;bcd0<=6; end
			3237: begin bcd3<=3;bcd2<=2;bcd1<=3;bcd0<=7; end
			3238: begin bcd3<=3;bcd2<=2;bcd1<=3;bcd0<=8; end
			3239: begin bcd3<=3;bcd2<=2;bcd1<=3;bcd0<=9; end
			3240: begin bcd3<=3;bcd2<=2;bcd1<=4;bcd0<=0; end
			3241: begin bcd3<=3;bcd2<=2;bcd1<=4;bcd0<=1; end
			3242: begin bcd3<=3;bcd2<=2;bcd1<=4;bcd0<=2; end
			3243: begin bcd3<=3;bcd2<=2;bcd1<=4;bcd0<=3; end
			3244: begin bcd3<=3;bcd2<=2;bcd1<=4;bcd0<=4; end
			3245: begin bcd3<=3;bcd2<=2;bcd1<=4;bcd0<=5; end
			3246: begin bcd3<=3;bcd2<=2;bcd1<=4;bcd0<=6; end
			3247: begin bcd3<=3;bcd2<=2;bcd1<=4;bcd0<=7; end
			3248: begin bcd3<=3;bcd2<=2;bcd1<=4;bcd0<=8; end
			3249: begin bcd3<=3;bcd2<=2;bcd1<=4;bcd0<=9; end
			3250: begin bcd3<=3;bcd2<=2;bcd1<=5;bcd0<=0; end
			3251: begin bcd3<=3;bcd2<=2;bcd1<=5;bcd0<=1; end
			3252: begin bcd3<=3;bcd2<=2;bcd1<=5;bcd0<=2; end
			3253: begin bcd3<=3;bcd2<=2;bcd1<=5;bcd0<=3; end
			3254: begin bcd3<=3;bcd2<=2;bcd1<=5;bcd0<=4; end
			3255: begin bcd3<=3;bcd2<=2;bcd1<=5;bcd0<=5; end
			3256: begin bcd3<=3;bcd2<=2;bcd1<=5;bcd0<=6; end
			3257: begin bcd3<=3;bcd2<=2;bcd1<=5;bcd0<=7; end
			3258: begin bcd3<=3;bcd2<=2;bcd1<=5;bcd0<=8; end
			3259: begin bcd3<=3;bcd2<=2;bcd1<=5;bcd0<=9; end
			3260: begin bcd3<=3;bcd2<=2;bcd1<=6;bcd0<=0; end
			3261: begin bcd3<=3;bcd2<=2;bcd1<=6;bcd0<=1; end
			3262: begin bcd3<=3;bcd2<=2;bcd1<=6;bcd0<=2; end
			3263: begin bcd3<=3;bcd2<=2;bcd1<=6;bcd0<=3; end
			3264: begin bcd3<=3;bcd2<=2;bcd1<=6;bcd0<=4; end
			3265: begin bcd3<=3;bcd2<=2;bcd1<=6;bcd0<=5; end
			3266: begin bcd3<=3;bcd2<=2;bcd1<=6;bcd0<=6; end
			3267: begin bcd3<=3;bcd2<=2;bcd1<=6;bcd0<=7; end
			3268: begin bcd3<=3;bcd2<=2;bcd1<=6;bcd0<=8; end
			3269: begin bcd3<=3;bcd2<=2;bcd1<=6;bcd0<=9; end
			3270: begin bcd3<=3;bcd2<=2;bcd1<=7;bcd0<=0; end
			3271: begin bcd3<=3;bcd2<=2;bcd1<=7;bcd0<=1; end
			3272: begin bcd3<=3;bcd2<=2;bcd1<=7;bcd0<=2; end
			3273: begin bcd3<=3;bcd2<=2;bcd1<=7;bcd0<=3; end
			3274: begin bcd3<=3;bcd2<=2;bcd1<=7;bcd0<=4; end
			3275: begin bcd3<=3;bcd2<=2;bcd1<=7;bcd0<=5; end
			3276: begin bcd3<=3;bcd2<=2;bcd1<=7;bcd0<=6; end
			3277: begin bcd3<=3;bcd2<=2;bcd1<=7;bcd0<=7; end
			3278: begin bcd3<=3;bcd2<=2;bcd1<=7;bcd0<=8; end
			3279: begin bcd3<=3;bcd2<=2;bcd1<=7;bcd0<=9; end
			3280: begin bcd3<=3;bcd2<=2;bcd1<=8;bcd0<=0; end
			3281: begin bcd3<=3;bcd2<=2;bcd1<=8;bcd0<=1; end
			3282: begin bcd3<=3;bcd2<=2;bcd1<=8;bcd0<=2; end
			3283: begin bcd3<=3;bcd2<=2;bcd1<=8;bcd0<=3; end
			3284: begin bcd3<=3;bcd2<=2;bcd1<=8;bcd0<=4; end
			3285: begin bcd3<=3;bcd2<=2;bcd1<=8;bcd0<=5; end
			3286: begin bcd3<=3;bcd2<=2;bcd1<=8;bcd0<=6; end
			3287: begin bcd3<=3;bcd2<=2;bcd1<=8;bcd0<=7; end
			3288: begin bcd3<=3;bcd2<=2;bcd1<=8;bcd0<=8; end
			3289: begin bcd3<=3;bcd2<=2;bcd1<=8;bcd0<=9; end
			3290: begin bcd3<=3;bcd2<=2;bcd1<=9;bcd0<=0; end
			3291: begin bcd3<=3;bcd2<=2;bcd1<=9;bcd0<=1; end
			3292: begin bcd3<=3;bcd2<=2;bcd1<=9;bcd0<=2; end
			3293: begin bcd3<=3;bcd2<=2;bcd1<=9;bcd0<=3; end
			3294: begin bcd3<=3;bcd2<=2;bcd1<=9;bcd0<=4; end
			3295: begin bcd3<=3;bcd2<=2;bcd1<=9;bcd0<=5; end
			3296: begin bcd3<=3;bcd2<=2;bcd1<=9;bcd0<=6; end
			3297: begin bcd3<=3;bcd2<=2;bcd1<=9;bcd0<=7; end
			3298: begin bcd3<=3;bcd2<=2;bcd1<=9;bcd0<=8; end
			3299: begin bcd3<=3;bcd2<=2;bcd1<=9;bcd0<=9; end
			3300: begin bcd3<=3;bcd2<=3;bcd1<=0;bcd0<=0; end
			3301: begin bcd3<=3;bcd2<=3;bcd1<=0;bcd0<=1; end
			3302: begin bcd3<=3;bcd2<=3;bcd1<=0;bcd0<=2; end
			3303: begin bcd3<=3;bcd2<=3;bcd1<=0;bcd0<=3; end
			3304: begin bcd3<=3;bcd2<=3;bcd1<=0;bcd0<=4; end
			3305: begin bcd3<=3;bcd2<=3;bcd1<=0;bcd0<=5; end
			3306: begin bcd3<=3;bcd2<=3;bcd1<=0;bcd0<=6; end
			3307: begin bcd3<=3;bcd2<=3;bcd1<=0;bcd0<=7; end
			3308: begin bcd3<=3;bcd2<=3;bcd1<=0;bcd0<=8; end
			3309: begin bcd3<=3;bcd2<=3;bcd1<=0;bcd0<=9; end
			3310: begin bcd3<=3;bcd2<=3;bcd1<=1;bcd0<=0; end
			3311: begin bcd3<=3;bcd2<=3;bcd1<=1;bcd0<=1; end
			3312: begin bcd3<=3;bcd2<=3;bcd1<=1;bcd0<=2; end
			3313: begin bcd3<=3;bcd2<=3;bcd1<=1;bcd0<=3; end
			3314: begin bcd3<=3;bcd2<=3;bcd1<=1;bcd0<=4; end
			3315: begin bcd3<=3;bcd2<=3;bcd1<=1;bcd0<=5; end
			3316: begin bcd3<=3;bcd2<=3;bcd1<=1;bcd0<=6; end
			3317: begin bcd3<=3;bcd2<=3;bcd1<=1;bcd0<=7; end
			3318: begin bcd3<=3;bcd2<=3;bcd1<=1;bcd0<=8; end
			3319: begin bcd3<=3;bcd2<=3;bcd1<=1;bcd0<=9; end
			3320: begin bcd3<=3;bcd2<=3;bcd1<=2;bcd0<=0; end
			3321: begin bcd3<=3;bcd2<=3;bcd1<=2;bcd0<=1; end
			3322: begin bcd3<=3;bcd2<=3;bcd1<=2;bcd0<=2; end
			3323: begin bcd3<=3;bcd2<=3;bcd1<=2;bcd0<=3; end
			3324: begin bcd3<=3;bcd2<=3;bcd1<=2;bcd0<=4; end
			3325: begin bcd3<=3;bcd2<=3;bcd1<=2;bcd0<=5; end
			3326: begin bcd3<=3;bcd2<=3;bcd1<=2;bcd0<=6; end
			3327: begin bcd3<=3;bcd2<=3;bcd1<=2;bcd0<=7; end
			3328: begin bcd3<=3;bcd2<=3;bcd1<=2;bcd0<=8; end
			3329: begin bcd3<=3;bcd2<=3;bcd1<=2;bcd0<=9; end
			3330: begin bcd3<=3;bcd2<=3;bcd1<=3;bcd0<=0; end
			3331: begin bcd3<=3;bcd2<=3;bcd1<=3;bcd0<=1; end
			3332: begin bcd3<=3;bcd2<=3;bcd1<=3;bcd0<=2; end
			3333: begin bcd3<=3;bcd2<=3;bcd1<=3;bcd0<=3; end
			3334: begin bcd3<=3;bcd2<=3;bcd1<=3;bcd0<=4; end
			3335: begin bcd3<=3;bcd2<=3;bcd1<=3;bcd0<=5; end
			3336: begin bcd3<=3;bcd2<=3;bcd1<=3;bcd0<=6; end
			3337: begin bcd3<=3;bcd2<=3;bcd1<=3;bcd0<=7; end
			3338: begin bcd3<=3;bcd2<=3;bcd1<=3;bcd0<=8; end
			3339: begin bcd3<=3;bcd2<=3;bcd1<=3;bcd0<=9; end
			3340: begin bcd3<=3;bcd2<=3;bcd1<=4;bcd0<=0; end
			3341: begin bcd3<=3;bcd2<=3;bcd1<=4;bcd0<=1; end
			3342: begin bcd3<=3;bcd2<=3;bcd1<=4;bcd0<=2; end
			3343: begin bcd3<=3;bcd2<=3;bcd1<=4;bcd0<=3; end
			3344: begin bcd3<=3;bcd2<=3;bcd1<=4;bcd0<=4; end
			3345: begin bcd3<=3;bcd2<=3;bcd1<=4;bcd0<=5; end
			3346: begin bcd3<=3;bcd2<=3;bcd1<=4;bcd0<=6; end
			3347: begin bcd3<=3;bcd2<=3;bcd1<=4;bcd0<=7; end
			3348: begin bcd3<=3;bcd2<=3;bcd1<=4;bcd0<=8; end
			3349: begin bcd3<=3;bcd2<=3;bcd1<=4;bcd0<=9; end
			3350: begin bcd3<=3;bcd2<=3;bcd1<=5;bcd0<=0; end
			3351: begin bcd3<=3;bcd2<=3;bcd1<=5;bcd0<=1; end
			3352: begin bcd3<=3;bcd2<=3;bcd1<=5;bcd0<=2; end
			3353: begin bcd3<=3;bcd2<=3;bcd1<=5;bcd0<=3; end
			3354: begin bcd3<=3;bcd2<=3;bcd1<=5;bcd0<=4; end
			3355: begin bcd3<=3;bcd2<=3;bcd1<=5;bcd0<=5; end
			3356: begin bcd3<=3;bcd2<=3;bcd1<=5;bcd0<=6; end
			3357: begin bcd3<=3;bcd2<=3;bcd1<=5;bcd0<=7; end
			3358: begin bcd3<=3;bcd2<=3;bcd1<=5;bcd0<=8; end
			3359: begin bcd3<=3;bcd2<=3;bcd1<=5;bcd0<=9; end
			3360: begin bcd3<=3;bcd2<=3;bcd1<=6;bcd0<=0; end
			3361: begin bcd3<=3;bcd2<=3;bcd1<=6;bcd0<=1; end
			3362: begin bcd3<=3;bcd2<=3;bcd1<=6;bcd0<=2; end
			3363: begin bcd3<=3;bcd2<=3;bcd1<=6;bcd0<=3; end
			3364: begin bcd3<=3;bcd2<=3;bcd1<=6;bcd0<=4; end
			3365: begin bcd3<=3;bcd2<=3;bcd1<=6;bcd0<=5; end
			3366: begin bcd3<=3;bcd2<=3;bcd1<=6;bcd0<=6; end
			3367: begin bcd3<=3;bcd2<=3;bcd1<=6;bcd0<=7; end
			3368: begin bcd3<=3;bcd2<=3;bcd1<=6;bcd0<=8; end
			3369: begin bcd3<=3;bcd2<=3;bcd1<=6;bcd0<=9; end
			3370: begin bcd3<=3;bcd2<=3;bcd1<=7;bcd0<=0; end
			3371: begin bcd3<=3;bcd2<=3;bcd1<=7;bcd0<=1; end
			3372: begin bcd3<=3;bcd2<=3;bcd1<=7;bcd0<=2; end
			3373: begin bcd3<=3;bcd2<=3;bcd1<=7;bcd0<=3; end
			3374: begin bcd3<=3;bcd2<=3;bcd1<=7;bcd0<=4; end
			3375: begin bcd3<=3;bcd2<=3;bcd1<=7;bcd0<=5; end
			3376: begin bcd3<=3;bcd2<=3;bcd1<=7;bcd0<=6; end
			3377: begin bcd3<=3;bcd2<=3;bcd1<=7;bcd0<=7; end
			3378: begin bcd3<=3;bcd2<=3;bcd1<=7;bcd0<=8; end
			3379: begin bcd3<=3;bcd2<=3;bcd1<=7;bcd0<=9; end
			3380: begin bcd3<=3;bcd2<=3;bcd1<=8;bcd0<=0; end
			3381: begin bcd3<=3;bcd2<=3;bcd1<=8;bcd0<=1; end
			3382: begin bcd3<=3;bcd2<=3;bcd1<=8;bcd0<=2; end
			3383: begin bcd3<=3;bcd2<=3;bcd1<=8;bcd0<=3; end
			3384: begin bcd3<=3;bcd2<=3;bcd1<=8;bcd0<=4; end
			3385: begin bcd3<=3;bcd2<=3;bcd1<=8;bcd0<=5; end
			3386: begin bcd3<=3;bcd2<=3;bcd1<=8;bcd0<=6; end
			3387: begin bcd3<=3;bcd2<=3;bcd1<=8;bcd0<=7; end
			3388: begin bcd3<=3;bcd2<=3;bcd1<=8;bcd0<=8; end
			3389: begin bcd3<=3;bcd2<=3;bcd1<=8;bcd0<=9; end
			3390: begin bcd3<=3;bcd2<=3;bcd1<=9;bcd0<=0; end
			3391: begin bcd3<=3;bcd2<=3;bcd1<=9;bcd0<=1; end
			3392: begin bcd3<=3;bcd2<=3;bcd1<=9;bcd0<=2; end
			3393: begin bcd3<=3;bcd2<=3;bcd1<=9;bcd0<=3; end
			3394: begin bcd3<=3;bcd2<=3;bcd1<=9;bcd0<=4; end
			3395: begin bcd3<=3;bcd2<=3;bcd1<=9;bcd0<=5; end
			3396: begin bcd3<=3;bcd2<=3;bcd1<=9;bcd0<=6; end
			3397: begin bcd3<=3;bcd2<=3;bcd1<=9;bcd0<=7; end
			3398: begin bcd3<=3;bcd2<=3;bcd1<=9;bcd0<=8; end
			3399: begin bcd3<=3;bcd2<=3;bcd1<=9;bcd0<=9; end
			3400: begin bcd3<=3;bcd2<=4;bcd1<=0;bcd0<=0; end
			3401: begin bcd3<=3;bcd2<=4;bcd1<=0;bcd0<=1; end
			3402: begin bcd3<=3;bcd2<=4;bcd1<=0;bcd0<=2; end
			3403: begin bcd3<=3;bcd2<=4;bcd1<=0;bcd0<=3; end
			3404: begin bcd3<=3;bcd2<=4;bcd1<=0;bcd0<=4; end
			3405: begin bcd3<=3;bcd2<=4;bcd1<=0;bcd0<=5; end
			3406: begin bcd3<=3;bcd2<=4;bcd1<=0;bcd0<=6; end
			3407: begin bcd3<=3;bcd2<=4;bcd1<=0;bcd0<=7; end
			3408: begin bcd3<=3;bcd2<=4;bcd1<=0;bcd0<=8; end
			3409: begin bcd3<=3;bcd2<=4;bcd1<=0;bcd0<=9; end
			3410: begin bcd3<=3;bcd2<=4;bcd1<=1;bcd0<=0; end
			3411: begin bcd3<=3;bcd2<=4;bcd1<=1;bcd0<=1; end
			3412: begin bcd3<=3;bcd2<=4;bcd1<=1;bcd0<=2; end
			3413: begin bcd3<=3;bcd2<=4;bcd1<=1;bcd0<=3; end
			3414: begin bcd3<=3;bcd2<=4;bcd1<=1;bcd0<=4; end
			3415: begin bcd3<=3;bcd2<=4;bcd1<=1;bcd0<=5; end
			3416: begin bcd3<=3;bcd2<=4;bcd1<=1;bcd0<=6; end
			3417: begin bcd3<=3;bcd2<=4;bcd1<=1;bcd0<=7; end
			3418: begin bcd3<=3;bcd2<=4;bcd1<=1;bcd0<=8; end
			3419: begin bcd3<=3;bcd2<=4;bcd1<=1;bcd0<=9; end
			3420: begin bcd3<=3;bcd2<=4;bcd1<=2;bcd0<=0; end
			3421: begin bcd3<=3;bcd2<=4;bcd1<=2;bcd0<=1; end
			3422: begin bcd3<=3;bcd2<=4;bcd1<=2;bcd0<=2; end
			3423: begin bcd3<=3;bcd2<=4;bcd1<=2;bcd0<=3; end
			3424: begin bcd3<=3;bcd2<=4;bcd1<=2;bcd0<=4; end
			3425: begin bcd3<=3;bcd2<=4;bcd1<=2;bcd0<=5; end
			3426: begin bcd3<=3;bcd2<=4;bcd1<=2;bcd0<=6; end
			3427: begin bcd3<=3;bcd2<=4;bcd1<=2;bcd0<=7; end
			3428: begin bcd3<=3;bcd2<=4;bcd1<=2;bcd0<=8; end
			3429: begin bcd3<=3;bcd2<=4;bcd1<=2;bcd0<=9; end
			3430: begin bcd3<=3;bcd2<=4;bcd1<=3;bcd0<=0; end
			3431: begin bcd3<=3;bcd2<=4;bcd1<=3;bcd0<=1; end
			3432: begin bcd3<=3;bcd2<=4;bcd1<=3;bcd0<=2; end
			3433: begin bcd3<=3;bcd2<=4;bcd1<=3;bcd0<=3; end
			3434: begin bcd3<=3;bcd2<=4;bcd1<=3;bcd0<=4; end
			3435: begin bcd3<=3;bcd2<=4;bcd1<=3;bcd0<=5; end
			3436: begin bcd3<=3;bcd2<=4;bcd1<=3;bcd0<=6; end
			3437: begin bcd3<=3;bcd2<=4;bcd1<=3;bcd0<=7; end
			3438: begin bcd3<=3;bcd2<=4;bcd1<=3;bcd0<=8; end
			3439: begin bcd3<=3;bcd2<=4;bcd1<=3;bcd0<=9; end
			3440: begin bcd3<=3;bcd2<=4;bcd1<=4;bcd0<=0; end
			3441: begin bcd3<=3;bcd2<=4;bcd1<=4;bcd0<=1; end
			3442: begin bcd3<=3;bcd2<=4;bcd1<=4;bcd0<=2; end
			3443: begin bcd3<=3;bcd2<=4;bcd1<=4;bcd0<=3; end
			3444: begin bcd3<=3;bcd2<=4;bcd1<=4;bcd0<=4; end
			3445: begin bcd3<=3;bcd2<=4;bcd1<=4;bcd0<=5; end
			3446: begin bcd3<=3;bcd2<=4;bcd1<=4;bcd0<=6; end
			3447: begin bcd3<=3;bcd2<=4;bcd1<=4;bcd0<=7; end
			3448: begin bcd3<=3;bcd2<=4;bcd1<=4;bcd0<=8; end
			3449: begin bcd3<=3;bcd2<=4;bcd1<=4;bcd0<=9; end
			3450: begin bcd3<=3;bcd2<=4;bcd1<=5;bcd0<=0; end
			3451: begin bcd3<=3;bcd2<=4;bcd1<=5;bcd0<=1; end
			3452: begin bcd3<=3;bcd2<=4;bcd1<=5;bcd0<=2; end
			3453: begin bcd3<=3;bcd2<=4;bcd1<=5;bcd0<=3; end
			3454: begin bcd3<=3;bcd2<=4;bcd1<=5;bcd0<=4; end
			3455: begin bcd3<=3;bcd2<=4;bcd1<=5;bcd0<=5; end
			3456: begin bcd3<=3;bcd2<=4;bcd1<=5;bcd0<=6; end
			3457: begin bcd3<=3;bcd2<=4;bcd1<=5;bcd0<=7; end
			3458: begin bcd3<=3;bcd2<=4;bcd1<=5;bcd0<=8; end
			3459: begin bcd3<=3;bcd2<=4;bcd1<=5;bcd0<=9; end
			3460: begin bcd3<=3;bcd2<=4;bcd1<=6;bcd0<=0; end
			3461: begin bcd3<=3;bcd2<=4;bcd1<=6;bcd0<=1; end
			3462: begin bcd3<=3;bcd2<=4;bcd1<=6;bcd0<=2; end
			3463: begin bcd3<=3;bcd2<=4;bcd1<=6;bcd0<=3; end
			3464: begin bcd3<=3;bcd2<=4;bcd1<=6;bcd0<=4; end
			3465: begin bcd3<=3;bcd2<=4;bcd1<=6;bcd0<=5; end
			3466: begin bcd3<=3;bcd2<=4;bcd1<=6;bcd0<=6; end
			3467: begin bcd3<=3;bcd2<=4;bcd1<=6;bcd0<=7; end
			3468: begin bcd3<=3;bcd2<=4;bcd1<=6;bcd0<=8; end
			3469: begin bcd3<=3;bcd2<=4;bcd1<=6;bcd0<=9; end
			3470: begin bcd3<=3;bcd2<=4;bcd1<=7;bcd0<=0; end
			3471: begin bcd3<=3;bcd2<=4;bcd1<=7;bcd0<=1; end
			3472: begin bcd3<=3;bcd2<=4;bcd1<=7;bcd0<=2; end
			3473: begin bcd3<=3;bcd2<=4;bcd1<=7;bcd0<=3; end
			3474: begin bcd3<=3;bcd2<=4;bcd1<=7;bcd0<=4; end
			3475: begin bcd3<=3;bcd2<=4;bcd1<=7;bcd0<=5; end
			3476: begin bcd3<=3;bcd2<=4;bcd1<=7;bcd0<=6; end
			3477: begin bcd3<=3;bcd2<=4;bcd1<=7;bcd0<=7; end
			3478: begin bcd3<=3;bcd2<=4;bcd1<=7;bcd0<=8; end
			3479: begin bcd3<=3;bcd2<=4;bcd1<=7;bcd0<=9; end
			3480: begin bcd3<=3;bcd2<=4;bcd1<=8;bcd0<=0; end
			3481: begin bcd3<=3;bcd2<=4;bcd1<=8;bcd0<=1; end
			3482: begin bcd3<=3;bcd2<=4;bcd1<=8;bcd0<=2; end
			3483: begin bcd3<=3;bcd2<=4;bcd1<=8;bcd0<=3; end
			3484: begin bcd3<=3;bcd2<=4;bcd1<=8;bcd0<=4; end
			3485: begin bcd3<=3;bcd2<=4;bcd1<=8;bcd0<=5; end
			3486: begin bcd3<=3;bcd2<=4;bcd1<=8;bcd0<=6; end
			3487: begin bcd3<=3;bcd2<=4;bcd1<=8;bcd0<=7; end
			3488: begin bcd3<=3;bcd2<=4;bcd1<=8;bcd0<=8; end
			3489: begin bcd3<=3;bcd2<=4;bcd1<=8;bcd0<=9; end
			3490: begin bcd3<=3;bcd2<=4;bcd1<=9;bcd0<=0; end
			3491: begin bcd3<=3;bcd2<=4;bcd1<=9;bcd0<=1; end
			3492: begin bcd3<=3;bcd2<=4;bcd1<=9;bcd0<=2; end
			3493: begin bcd3<=3;bcd2<=4;bcd1<=9;bcd0<=3; end
			3494: begin bcd3<=3;bcd2<=4;bcd1<=9;bcd0<=4; end
			3495: begin bcd3<=3;bcd2<=4;bcd1<=9;bcd0<=5; end
			3496: begin bcd3<=3;bcd2<=4;bcd1<=9;bcd0<=6; end
			3497: begin bcd3<=3;bcd2<=4;bcd1<=9;bcd0<=7; end
			3498: begin bcd3<=3;bcd2<=4;bcd1<=9;bcd0<=8; end
			3499: begin bcd3<=3;bcd2<=4;bcd1<=9;bcd0<=9; end
			3500: begin bcd3<=3;bcd2<=5;bcd1<=0;bcd0<=0; end
			3501: begin bcd3<=3;bcd2<=5;bcd1<=0;bcd0<=1; end
			3502: begin bcd3<=3;bcd2<=5;bcd1<=0;bcd0<=2; end
			3503: begin bcd3<=3;bcd2<=5;bcd1<=0;bcd0<=3; end
			3504: begin bcd3<=3;bcd2<=5;bcd1<=0;bcd0<=4; end
			3505: begin bcd3<=3;bcd2<=5;bcd1<=0;bcd0<=5; end
			3506: begin bcd3<=3;bcd2<=5;bcd1<=0;bcd0<=6; end
			3507: begin bcd3<=3;bcd2<=5;bcd1<=0;bcd0<=7; end
			3508: begin bcd3<=3;bcd2<=5;bcd1<=0;bcd0<=8; end
			3509: begin bcd3<=3;bcd2<=5;bcd1<=0;bcd0<=9; end
			3510: begin bcd3<=3;bcd2<=5;bcd1<=1;bcd0<=0; end
			3511: begin bcd3<=3;bcd2<=5;bcd1<=1;bcd0<=1; end
			3512: begin bcd3<=3;bcd2<=5;bcd1<=1;bcd0<=2; end
			3513: begin bcd3<=3;bcd2<=5;bcd1<=1;bcd0<=3; end
			3514: begin bcd3<=3;bcd2<=5;bcd1<=1;bcd0<=4; end
			3515: begin bcd3<=3;bcd2<=5;bcd1<=1;bcd0<=5; end
			3516: begin bcd3<=3;bcd2<=5;bcd1<=1;bcd0<=6; end
			3517: begin bcd3<=3;bcd2<=5;bcd1<=1;bcd0<=7; end
			3518: begin bcd3<=3;bcd2<=5;bcd1<=1;bcd0<=8; end
			3519: begin bcd3<=3;bcd2<=5;bcd1<=1;bcd0<=9; end
			3520: begin bcd3<=3;bcd2<=5;bcd1<=2;bcd0<=0; end
			3521: begin bcd3<=3;bcd2<=5;bcd1<=2;bcd0<=1; end
			3522: begin bcd3<=3;bcd2<=5;bcd1<=2;bcd0<=2; end
			3523: begin bcd3<=3;bcd2<=5;bcd1<=2;bcd0<=3; end
			3524: begin bcd3<=3;bcd2<=5;bcd1<=2;bcd0<=4; end
			3525: begin bcd3<=3;bcd2<=5;bcd1<=2;bcd0<=5; end
			3526: begin bcd3<=3;bcd2<=5;bcd1<=2;bcd0<=6; end
			3527: begin bcd3<=3;bcd2<=5;bcd1<=2;bcd0<=7; end
			3528: begin bcd3<=3;bcd2<=5;bcd1<=2;bcd0<=8; end
			3529: begin bcd3<=3;bcd2<=5;bcd1<=2;bcd0<=9; end
			3530: begin bcd3<=3;bcd2<=5;bcd1<=3;bcd0<=0; end
			3531: begin bcd3<=3;bcd2<=5;bcd1<=3;bcd0<=1; end
			3532: begin bcd3<=3;bcd2<=5;bcd1<=3;bcd0<=2; end
			3533: begin bcd3<=3;bcd2<=5;bcd1<=3;bcd0<=3; end
			3534: begin bcd3<=3;bcd2<=5;bcd1<=3;bcd0<=4; end
			3535: begin bcd3<=3;bcd2<=5;bcd1<=3;bcd0<=5; end
			3536: begin bcd3<=3;bcd2<=5;bcd1<=3;bcd0<=6; end
			3537: begin bcd3<=3;bcd2<=5;bcd1<=3;bcd0<=7; end
			3538: begin bcd3<=3;bcd2<=5;bcd1<=3;bcd0<=8; end
			3539: begin bcd3<=3;bcd2<=5;bcd1<=3;bcd0<=9; end
			3540: begin bcd3<=3;bcd2<=5;bcd1<=4;bcd0<=0; end
			3541: begin bcd3<=3;bcd2<=5;bcd1<=4;bcd0<=1; end
			3542: begin bcd3<=3;bcd2<=5;bcd1<=4;bcd0<=2; end
			3543: begin bcd3<=3;bcd2<=5;bcd1<=4;bcd0<=3; end
			3544: begin bcd3<=3;bcd2<=5;bcd1<=4;bcd0<=4; end
			3545: begin bcd3<=3;bcd2<=5;bcd1<=4;bcd0<=5; end
			3546: begin bcd3<=3;bcd2<=5;bcd1<=4;bcd0<=6; end
			3547: begin bcd3<=3;bcd2<=5;bcd1<=4;bcd0<=7; end
			3548: begin bcd3<=3;bcd2<=5;bcd1<=4;bcd0<=8; end
			3549: begin bcd3<=3;bcd2<=5;bcd1<=4;bcd0<=9; end
			3550: begin bcd3<=3;bcd2<=5;bcd1<=5;bcd0<=0; end
			3551: begin bcd3<=3;bcd2<=5;bcd1<=5;bcd0<=1; end
			3552: begin bcd3<=3;bcd2<=5;bcd1<=5;bcd0<=2; end
			3553: begin bcd3<=3;bcd2<=5;bcd1<=5;bcd0<=3; end
			3554: begin bcd3<=3;bcd2<=5;bcd1<=5;bcd0<=4; end
			3555: begin bcd3<=3;bcd2<=5;bcd1<=5;bcd0<=5; end
			3556: begin bcd3<=3;bcd2<=5;bcd1<=5;bcd0<=6; end
			3557: begin bcd3<=3;bcd2<=5;bcd1<=5;bcd0<=7; end
			3558: begin bcd3<=3;bcd2<=5;bcd1<=5;bcd0<=8; end
			3559: begin bcd3<=3;bcd2<=5;bcd1<=5;bcd0<=9; end
			3560: begin bcd3<=3;bcd2<=5;bcd1<=6;bcd0<=0; end
			3561: begin bcd3<=3;bcd2<=5;bcd1<=6;bcd0<=1; end
			3562: begin bcd3<=3;bcd2<=5;bcd1<=6;bcd0<=2; end
			3563: begin bcd3<=3;bcd2<=5;bcd1<=6;bcd0<=3; end
			3564: begin bcd3<=3;bcd2<=5;bcd1<=6;bcd0<=4; end
			3565: begin bcd3<=3;bcd2<=5;bcd1<=6;bcd0<=5; end
			3566: begin bcd3<=3;bcd2<=5;bcd1<=6;bcd0<=6; end
			3567: begin bcd3<=3;bcd2<=5;bcd1<=6;bcd0<=7; end
			3568: begin bcd3<=3;bcd2<=5;bcd1<=6;bcd0<=8; end
			3569: begin bcd3<=3;bcd2<=5;bcd1<=6;bcd0<=9; end
			3570: begin bcd3<=3;bcd2<=5;bcd1<=7;bcd0<=0; end
			3571: begin bcd3<=3;bcd2<=5;bcd1<=7;bcd0<=1; end
			3572: begin bcd3<=3;bcd2<=5;bcd1<=7;bcd0<=2; end
			3573: begin bcd3<=3;bcd2<=5;bcd1<=7;bcd0<=3; end
			3574: begin bcd3<=3;bcd2<=5;bcd1<=7;bcd0<=4; end
			3575: begin bcd3<=3;bcd2<=5;bcd1<=7;bcd0<=5; end
			3576: begin bcd3<=3;bcd2<=5;bcd1<=7;bcd0<=6; end
			3577: begin bcd3<=3;bcd2<=5;bcd1<=7;bcd0<=7; end
			3578: begin bcd3<=3;bcd2<=5;bcd1<=7;bcd0<=8; end
			3579: begin bcd3<=3;bcd2<=5;bcd1<=7;bcd0<=9; end
			3580: begin bcd3<=3;bcd2<=5;bcd1<=8;bcd0<=0; end
			3581: begin bcd3<=3;bcd2<=5;bcd1<=8;bcd0<=1; end
			3582: begin bcd3<=3;bcd2<=5;bcd1<=8;bcd0<=2; end
			3583: begin bcd3<=3;bcd2<=5;bcd1<=8;bcd0<=3; end
			3584: begin bcd3<=3;bcd2<=5;bcd1<=8;bcd0<=4; end
			3585: begin bcd3<=3;bcd2<=5;bcd1<=8;bcd0<=5; end
			3586: begin bcd3<=3;bcd2<=5;bcd1<=8;bcd0<=6; end
			3587: begin bcd3<=3;bcd2<=5;bcd1<=8;bcd0<=7; end
			3588: begin bcd3<=3;bcd2<=5;bcd1<=8;bcd0<=8; end
			3589: begin bcd3<=3;bcd2<=5;bcd1<=8;bcd0<=9; end
			3590: begin bcd3<=3;bcd2<=5;bcd1<=9;bcd0<=0; end
			3591: begin bcd3<=3;bcd2<=5;bcd1<=9;bcd0<=1; end
			3592: begin bcd3<=3;bcd2<=5;bcd1<=9;bcd0<=2; end
			3593: begin bcd3<=3;bcd2<=5;bcd1<=9;bcd0<=3; end
			3594: begin bcd3<=3;bcd2<=5;bcd1<=9;bcd0<=4; end
			3595: begin bcd3<=3;bcd2<=5;bcd1<=9;bcd0<=5; end
			3596: begin bcd3<=3;bcd2<=5;bcd1<=9;bcd0<=6; end
			3597: begin bcd3<=3;bcd2<=5;bcd1<=9;bcd0<=7; end
			3598: begin bcd3<=3;bcd2<=5;bcd1<=9;bcd0<=8; end
			3599: begin bcd3<=3;bcd2<=5;bcd1<=9;bcd0<=9; end
			3600: begin bcd3<=3;bcd2<=6;bcd1<=0;bcd0<=0; end
			3601: begin bcd3<=3;bcd2<=6;bcd1<=0;bcd0<=1; end
			3602: begin bcd3<=3;bcd2<=6;bcd1<=0;bcd0<=2; end
			3603: begin bcd3<=3;bcd2<=6;bcd1<=0;bcd0<=3; end
			3604: begin bcd3<=3;bcd2<=6;bcd1<=0;bcd0<=4; end
			3605: begin bcd3<=3;bcd2<=6;bcd1<=0;bcd0<=5; end
			3606: begin bcd3<=3;bcd2<=6;bcd1<=0;bcd0<=6; end
			3607: begin bcd3<=3;bcd2<=6;bcd1<=0;bcd0<=7; end
			3608: begin bcd3<=3;bcd2<=6;bcd1<=0;bcd0<=8; end
			3609: begin bcd3<=3;bcd2<=6;bcd1<=0;bcd0<=9; end
			3610: begin bcd3<=3;bcd2<=6;bcd1<=1;bcd0<=0; end
			3611: begin bcd3<=3;bcd2<=6;bcd1<=1;bcd0<=1; end
			3612: begin bcd3<=3;bcd2<=6;bcd1<=1;bcd0<=2; end
			3613: begin bcd3<=3;bcd2<=6;bcd1<=1;bcd0<=3; end
			3614: begin bcd3<=3;bcd2<=6;bcd1<=1;bcd0<=4; end
			3615: begin bcd3<=3;bcd2<=6;bcd1<=1;bcd0<=5; end
			3616: begin bcd3<=3;bcd2<=6;bcd1<=1;bcd0<=6; end
			3617: begin bcd3<=3;bcd2<=6;bcd1<=1;bcd0<=7; end
			3618: begin bcd3<=3;bcd2<=6;bcd1<=1;bcd0<=8; end
			3619: begin bcd3<=3;bcd2<=6;bcd1<=1;bcd0<=9; end
			3620: begin bcd3<=3;bcd2<=6;bcd1<=2;bcd0<=0; end
			3621: begin bcd3<=3;bcd2<=6;bcd1<=2;bcd0<=1; end
			3622: begin bcd3<=3;bcd2<=6;bcd1<=2;bcd0<=2; end
			3623: begin bcd3<=3;bcd2<=6;bcd1<=2;bcd0<=3; end
			3624: begin bcd3<=3;bcd2<=6;bcd1<=2;bcd0<=4; end
			3625: begin bcd3<=3;bcd2<=6;bcd1<=2;bcd0<=5; end
			3626: begin bcd3<=3;bcd2<=6;bcd1<=2;bcd0<=6; end
			3627: begin bcd3<=3;bcd2<=6;bcd1<=2;bcd0<=7; end
			3628: begin bcd3<=3;bcd2<=6;bcd1<=2;bcd0<=8; end
			3629: begin bcd3<=3;bcd2<=6;bcd1<=2;bcd0<=9; end
			3630: begin bcd3<=3;bcd2<=6;bcd1<=3;bcd0<=0; end
			3631: begin bcd3<=3;bcd2<=6;bcd1<=3;bcd0<=1; end
			3632: begin bcd3<=3;bcd2<=6;bcd1<=3;bcd0<=2; end
			3633: begin bcd3<=3;bcd2<=6;bcd1<=3;bcd0<=3; end
			3634: begin bcd3<=3;bcd2<=6;bcd1<=3;bcd0<=4; end
			3635: begin bcd3<=3;bcd2<=6;bcd1<=3;bcd0<=5; end
			3636: begin bcd3<=3;bcd2<=6;bcd1<=3;bcd0<=6; end
			3637: begin bcd3<=3;bcd2<=6;bcd1<=3;bcd0<=7; end
			3638: begin bcd3<=3;bcd2<=6;bcd1<=3;bcd0<=8; end
			3639: begin bcd3<=3;bcd2<=6;bcd1<=3;bcd0<=9; end
			3640: begin bcd3<=3;bcd2<=6;bcd1<=4;bcd0<=0; end
			3641: begin bcd3<=3;bcd2<=6;bcd1<=4;bcd0<=1; end
			3642: begin bcd3<=3;bcd2<=6;bcd1<=4;bcd0<=2; end
			3643: begin bcd3<=3;bcd2<=6;bcd1<=4;bcd0<=3; end
			3644: begin bcd3<=3;bcd2<=6;bcd1<=4;bcd0<=4; end
			3645: begin bcd3<=3;bcd2<=6;bcd1<=4;bcd0<=5; end
			3646: begin bcd3<=3;bcd2<=6;bcd1<=4;bcd0<=6; end
			3647: begin bcd3<=3;bcd2<=6;bcd1<=4;bcd0<=7; end
			3648: begin bcd3<=3;bcd2<=6;bcd1<=4;bcd0<=8; end
			3649: begin bcd3<=3;bcd2<=6;bcd1<=4;bcd0<=9; end
			3650: begin bcd3<=3;bcd2<=6;bcd1<=5;bcd0<=0; end
			3651: begin bcd3<=3;bcd2<=6;bcd1<=5;bcd0<=1; end
			3652: begin bcd3<=3;bcd2<=6;bcd1<=5;bcd0<=2; end
			3653: begin bcd3<=3;bcd2<=6;bcd1<=5;bcd0<=3; end
			3654: begin bcd3<=3;bcd2<=6;bcd1<=5;bcd0<=4; end
			3655: begin bcd3<=3;bcd2<=6;bcd1<=5;bcd0<=5; end
			3656: begin bcd3<=3;bcd2<=6;bcd1<=5;bcd0<=6; end
			3657: begin bcd3<=3;bcd2<=6;bcd1<=5;bcd0<=7; end
			3658: begin bcd3<=3;bcd2<=6;bcd1<=5;bcd0<=8; end
			3659: begin bcd3<=3;bcd2<=6;bcd1<=5;bcd0<=9; end
			3660: begin bcd3<=3;bcd2<=6;bcd1<=6;bcd0<=0; end
			3661: begin bcd3<=3;bcd2<=6;bcd1<=6;bcd0<=1; end
			3662: begin bcd3<=3;bcd2<=6;bcd1<=6;bcd0<=2; end
			3663: begin bcd3<=3;bcd2<=6;bcd1<=6;bcd0<=3; end
			3664: begin bcd3<=3;bcd2<=6;bcd1<=6;bcd0<=4; end
			3665: begin bcd3<=3;bcd2<=6;bcd1<=6;bcd0<=5; end
			3666: begin bcd3<=3;bcd2<=6;bcd1<=6;bcd0<=6; end
			3667: begin bcd3<=3;bcd2<=6;bcd1<=6;bcd0<=7; end
			3668: begin bcd3<=3;bcd2<=6;bcd1<=6;bcd0<=8; end
			3669: begin bcd3<=3;bcd2<=6;bcd1<=6;bcd0<=9; end
			3670: begin bcd3<=3;bcd2<=6;bcd1<=7;bcd0<=0; end
			3671: begin bcd3<=3;bcd2<=6;bcd1<=7;bcd0<=1; end
			3672: begin bcd3<=3;bcd2<=6;bcd1<=7;bcd0<=2; end
			3673: begin bcd3<=3;bcd2<=6;bcd1<=7;bcd0<=3; end
			3674: begin bcd3<=3;bcd2<=6;bcd1<=7;bcd0<=4; end
			3675: begin bcd3<=3;bcd2<=6;bcd1<=7;bcd0<=5; end
			3676: begin bcd3<=3;bcd2<=6;bcd1<=7;bcd0<=6; end
			3677: begin bcd3<=3;bcd2<=6;bcd1<=7;bcd0<=7; end
			3678: begin bcd3<=3;bcd2<=6;bcd1<=7;bcd0<=8; end
			3679: begin bcd3<=3;bcd2<=6;bcd1<=7;bcd0<=9; end
			3680: begin bcd3<=3;bcd2<=6;bcd1<=8;bcd0<=0; end
			3681: begin bcd3<=3;bcd2<=6;bcd1<=8;bcd0<=1; end
			3682: begin bcd3<=3;bcd2<=6;bcd1<=8;bcd0<=2; end
			3683: begin bcd3<=3;bcd2<=6;bcd1<=8;bcd0<=3; end
			3684: begin bcd3<=3;bcd2<=6;bcd1<=8;bcd0<=4; end
			3685: begin bcd3<=3;bcd2<=6;bcd1<=8;bcd0<=5; end
			3686: begin bcd3<=3;bcd2<=6;bcd1<=8;bcd0<=6; end
			3687: begin bcd3<=3;bcd2<=6;bcd1<=8;bcd0<=7; end
			3688: begin bcd3<=3;bcd2<=6;bcd1<=8;bcd0<=8; end
			3689: begin bcd3<=3;bcd2<=6;bcd1<=8;bcd0<=9; end
			3690: begin bcd3<=3;bcd2<=6;bcd1<=9;bcd0<=0; end
			3691: begin bcd3<=3;bcd2<=6;bcd1<=9;bcd0<=1; end
			3692: begin bcd3<=3;bcd2<=6;bcd1<=9;bcd0<=2; end
			3693: begin bcd3<=3;bcd2<=6;bcd1<=9;bcd0<=3; end
			3694: begin bcd3<=3;bcd2<=6;bcd1<=9;bcd0<=4; end
			3695: begin bcd3<=3;bcd2<=6;bcd1<=9;bcd0<=5; end
			3696: begin bcd3<=3;bcd2<=6;bcd1<=9;bcd0<=6; end
			3697: begin bcd3<=3;bcd2<=6;bcd1<=9;bcd0<=7; end
			3698: begin bcd3<=3;bcd2<=6;bcd1<=9;bcd0<=8; end
			3699: begin bcd3<=3;bcd2<=6;bcd1<=9;bcd0<=9; end
			3700: begin bcd3<=3;bcd2<=7;bcd1<=0;bcd0<=0; end
			3701: begin bcd3<=3;bcd2<=7;bcd1<=0;bcd0<=1; end
			3702: begin bcd3<=3;bcd2<=7;bcd1<=0;bcd0<=2; end
			3703: begin bcd3<=3;bcd2<=7;bcd1<=0;bcd0<=3; end
			3704: begin bcd3<=3;bcd2<=7;bcd1<=0;bcd0<=4; end
			3705: begin bcd3<=3;bcd2<=7;bcd1<=0;bcd0<=5; end
			3706: begin bcd3<=3;bcd2<=7;bcd1<=0;bcd0<=6; end
			3707: begin bcd3<=3;bcd2<=7;bcd1<=0;bcd0<=7; end
			3708: begin bcd3<=3;bcd2<=7;bcd1<=0;bcd0<=8; end
			3709: begin bcd3<=3;bcd2<=7;bcd1<=0;bcd0<=9; end
			3710: begin bcd3<=3;bcd2<=7;bcd1<=1;bcd0<=0; end
			3711: begin bcd3<=3;bcd2<=7;bcd1<=1;bcd0<=1; end
			3712: begin bcd3<=3;bcd2<=7;bcd1<=1;bcd0<=2; end
			3713: begin bcd3<=3;bcd2<=7;bcd1<=1;bcd0<=3; end
			3714: begin bcd3<=3;bcd2<=7;bcd1<=1;bcd0<=4; end
			3715: begin bcd3<=3;bcd2<=7;bcd1<=1;bcd0<=5; end
			3716: begin bcd3<=3;bcd2<=7;bcd1<=1;bcd0<=6; end
			3717: begin bcd3<=3;bcd2<=7;bcd1<=1;bcd0<=7; end
			3718: begin bcd3<=3;bcd2<=7;bcd1<=1;bcd0<=8; end
			3719: begin bcd3<=3;bcd2<=7;bcd1<=1;bcd0<=9; end
			3720: begin bcd3<=3;bcd2<=7;bcd1<=2;bcd0<=0; end
			3721: begin bcd3<=3;bcd2<=7;bcd1<=2;bcd0<=1; end
			3722: begin bcd3<=3;bcd2<=7;bcd1<=2;bcd0<=2; end
			3723: begin bcd3<=3;bcd2<=7;bcd1<=2;bcd0<=3; end
			3724: begin bcd3<=3;bcd2<=7;bcd1<=2;bcd0<=4; end
			3725: begin bcd3<=3;bcd2<=7;bcd1<=2;bcd0<=5; end
			3726: begin bcd3<=3;bcd2<=7;bcd1<=2;bcd0<=6; end
			3727: begin bcd3<=3;bcd2<=7;bcd1<=2;bcd0<=7; end
			3728: begin bcd3<=3;bcd2<=7;bcd1<=2;bcd0<=8; end
			3729: begin bcd3<=3;bcd2<=7;bcd1<=2;bcd0<=9; end
			3730: begin bcd3<=3;bcd2<=7;bcd1<=3;bcd0<=0; end
			3731: begin bcd3<=3;bcd2<=7;bcd1<=3;bcd0<=1; end
			3732: begin bcd3<=3;bcd2<=7;bcd1<=3;bcd0<=2; end
			3733: begin bcd3<=3;bcd2<=7;bcd1<=3;bcd0<=3; end
			3734: begin bcd3<=3;bcd2<=7;bcd1<=3;bcd0<=4; end
			3735: begin bcd3<=3;bcd2<=7;bcd1<=3;bcd0<=5; end
			3736: begin bcd3<=3;bcd2<=7;bcd1<=3;bcd0<=6; end
			3737: begin bcd3<=3;bcd2<=7;bcd1<=3;bcd0<=7; end
			3738: begin bcd3<=3;bcd2<=7;bcd1<=3;bcd0<=8; end
			3739: begin bcd3<=3;bcd2<=7;bcd1<=3;bcd0<=9; end
			3740: begin bcd3<=3;bcd2<=7;bcd1<=4;bcd0<=0; end
			3741: begin bcd3<=3;bcd2<=7;bcd1<=4;bcd0<=1; end
			3742: begin bcd3<=3;bcd2<=7;bcd1<=4;bcd0<=2; end
			3743: begin bcd3<=3;bcd2<=7;bcd1<=4;bcd0<=3; end
			3744: begin bcd3<=3;bcd2<=7;bcd1<=4;bcd0<=4; end
			3745: begin bcd3<=3;bcd2<=7;bcd1<=4;bcd0<=5; end
			3746: begin bcd3<=3;bcd2<=7;bcd1<=4;bcd0<=6; end
			3747: begin bcd3<=3;bcd2<=7;bcd1<=4;bcd0<=7; end
			3748: begin bcd3<=3;bcd2<=7;bcd1<=4;bcd0<=8; end
			3749: begin bcd3<=3;bcd2<=7;bcd1<=4;bcd0<=9; end
			3750: begin bcd3<=3;bcd2<=7;bcd1<=5;bcd0<=0; end
			3751: begin bcd3<=3;bcd2<=7;bcd1<=5;bcd0<=1; end
			3752: begin bcd3<=3;bcd2<=7;bcd1<=5;bcd0<=2; end
			3753: begin bcd3<=3;bcd2<=7;bcd1<=5;bcd0<=3; end
			3754: begin bcd3<=3;bcd2<=7;bcd1<=5;bcd0<=4; end
			3755: begin bcd3<=3;bcd2<=7;bcd1<=5;bcd0<=5; end
			3756: begin bcd3<=3;bcd2<=7;bcd1<=5;bcd0<=6; end
			3757: begin bcd3<=3;bcd2<=7;bcd1<=5;bcd0<=7; end
			3758: begin bcd3<=3;bcd2<=7;bcd1<=5;bcd0<=8; end
			3759: begin bcd3<=3;bcd2<=7;bcd1<=5;bcd0<=9; end
			3760: begin bcd3<=3;bcd2<=7;bcd1<=6;bcd0<=0; end
			3761: begin bcd3<=3;bcd2<=7;bcd1<=6;bcd0<=1; end
			3762: begin bcd3<=3;bcd2<=7;bcd1<=6;bcd0<=2; end
			3763: begin bcd3<=3;bcd2<=7;bcd1<=6;bcd0<=3; end
			3764: begin bcd3<=3;bcd2<=7;bcd1<=6;bcd0<=4; end
			3765: begin bcd3<=3;bcd2<=7;bcd1<=6;bcd0<=5; end
			3766: begin bcd3<=3;bcd2<=7;bcd1<=6;bcd0<=6; end
			3767: begin bcd3<=3;bcd2<=7;bcd1<=6;bcd0<=7; end
			3768: begin bcd3<=3;bcd2<=7;bcd1<=6;bcd0<=8; end
			3769: begin bcd3<=3;bcd2<=7;bcd1<=6;bcd0<=9; end
			3770: begin bcd3<=3;bcd2<=7;bcd1<=7;bcd0<=0; end
			3771: begin bcd3<=3;bcd2<=7;bcd1<=7;bcd0<=1; end
			3772: begin bcd3<=3;bcd2<=7;bcd1<=7;bcd0<=2; end
			3773: begin bcd3<=3;bcd2<=7;bcd1<=7;bcd0<=3; end
			3774: begin bcd3<=3;bcd2<=7;bcd1<=7;bcd0<=4; end
			3775: begin bcd3<=3;bcd2<=7;bcd1<=7;bcd0<=5; end
			3776: begin bcd3<=3;bcd2<=7;bcd1<=7;bcd0<=6; end
			3777: begin bcd3<=3;bcd2<=7;bcd1<=7;bcd0<=7; end
			3778: begin bcd3<=3;bcd2<=7;bcd1<=7;bcd0<=8; end
			3779: begin bcd3<=3;bcd2<=7;bcd1<=7;bcd0<=9; end
			3780: begin bcd3<=3;bcd2<=7;bcd1<=8;bcd0<=0; end
			3781: begin bcd3<=3;bcd2<=7;bcd1<=8;bcd0<=1; end
			3782: begin bcd3<=3;bcd2<=7;bcd1<=8;bcd0<=2; end
			3783: begin bcd3<=3;bcd2<=7;bcd1<=8;bcd0<=3; end
			3784: begin bcd3<=3;bcd2<=7;bcd1<=8;bcd0<=4; end
			3785: begin bcd3<=3;bcd2<=7;bcd1<=8;bcd0<=5; end
			3786: begin bcd3<=3;bcd2<=7;bcd1<=8;bcd0<=6; end
			3787: begin bcd3<=3;bcd2<=7;bcd1<=8;bcd0<=7; end
			3788: begin bcd3<=3;bcd2<=7;bcd1<=8;bcd0<=8; end
			3789: begin bcd3<=3;bcd2<=7;bcd1<=8;bcd0<=9; end
			3790: begin bcd3<=3;bcd2<=7;bcd1<=9;bcd0<=0; end
			3791: begin bcd3<=3;bcd2<=7;bcd1<=9;bcd0<=1; end
			3792: begin bcd3<=3;bcd2<=7;bcd1<=9;bcd0<=2; end
			3793: begin bcd3<=3;bcd2<=7;bcd1<=9;bcd0<=3; end
			3794: begin bcd3<=3;bcd2<=7;bcd1<=9;bcd0<=4; end
			3795: begin bcd3<=3;bcd2<=7;bcd1<=9;bcd0<=5; end
			3796: begin bcd3<=3;bcd2<=7;bcd1<=9;bcd0<=6; end
			3797: begin bcd3<=3;bcd2<=7;bcd1<=9;bcd0<=7; end
			3798: begin bcd3<=3;bcd2<=7;bcd1<=9;bcd0<=8; end
			3799: begin bcd3<=3;bcd2<=7;bcd1<=9;bcd0<=9; end
			3800: begin bcd3<=3;bcd2<=8;bcd1<=0;bcd0<=0; end
			3801: begin bcd3<=3;bcd2<=8;bcd1<=0;bcd0<=1; end
			3802: begin bcd3<=3;bcd2<=8;bcd1<=0;bcd0<=2; end
			3803: begin bcd3<=3;bcd2<=8;bcd1<=0;bcd0<=3; end
			3804: begin bcd3<=3;bcd2<=8;bcd1<=0;bcd0<=4; end
			3805: begin bcd3<=3;bcd2<=8;bcd1<=0;bcd0<=5; end
			3806: begin bcd3<=3;bcd2<=8;bcd1<=0;bcd0<=6; end
			3807: begin bcd3<=3;bcd2<=8;bcd1<=0;bcd0<=7; end
			3808: begin bcd3<=3;bcd2<=8;bcd1<=0;bcd0<=8; end
			3809: begin bcd3<=3;bcd2<=8;bcd1<=0;bcd0<=9; end
			3810: begin bcd3<=3;bcd2<=8;bcd1<=1;bcd0<=0; end
			3811: begin bcd3<=3;bcd2<=8;bcd1<=1;bcd0<=1; end
			3812: begin bcd3<=3;bcd2<=8;bcd1<=1;bcd0<=2; end
			3813: begin bcd3<=3;bcd2<=8;bcd1<=1;bcd0<=3; end
			3814: begin bcd3<=3;bcd2<=8;bcd1<=1;bcd0<=4; end
			3815: begin bcd3<=3;bcd2<=8;bcd1<=1;bcd0<=5; end
			3816: begin bcd3<=3;bcd2<=8;bcd1<=1;bcd0<=6; end
			3817: begin bcd3<=3;bcd2<=8;bcd1<=1;bcd0<=7; end
			3818: begin bcd3<=3;bcd2<=8;bcd1<=1;bcd0<=8; end
			3819: begin bcd3<=3;bcd2<=8;bcd1<=1;bcd0<=9; end
			3820: begin bcd3<=3;bcd2<=8;bcd1<=2;bcd0<=0; end
			3821: begin bcd3<=3;bcd2<=8;bcd1<=2;bcd0<=1; end
			3822: begin bcd3<=3;bcd2<=8;bcd1<=2;bcd0<=2; end
			3823: begin bcd3<=3;bcd2<=8;bcd1<=2;bcd0<=3; end
			3824: begin bcd3<=3;bcd2<=8;bcd1<=2;bcd0<=4; end
			3825: begin bcd3<=3;bcd2<=8;bcd1<=2;bcd0<=5; end
			3826: begin bcd3<=3;bcd2<=8;bcd1<=2;bcd0<=6; end
			3827: begin bcd3<=3;bcd2<=8;bcd1<=2;bcd0<=7; end
			3828: begin bcd3<=3;bcd2<=8;bcd1<=2;bcd0<=8; end
			3829: begin bcd3<=3;bcd2<=8;bcd1<=2;bcd0<=9; end
			3830: begin bcd3<=3;bcd2<=8;bcd1<=3;bcd0<=0; end
			3831: begin bcd3<=3;bcd2<=8;bcd1<=3;bcd0<=1; end
			3832: begin bcd3<=3;bcd2<=8;bcd1<=3;bcd0<=2; end
			3833: begin bcd3<=3;bcd2<=8;bcd1<=3;bcd0<=3; end
			3834: begin bcd3<=3;bcd2<=8;bcd1<=3;bcd0<=4; end
			3835: begin bcd3<=3;bcd2<=8;bcd1<=3;bcd0<=5; end
			3836: begin bcd3<=3;bcd2<=8;bcd1<=3;bcd0<=6; end
			3837: begin bcd3<=3;bcd2<=8;bcd1<=3;bcd0<=7; end
			3838: begin bcd3<=3;bcd2<=8;bcd1<=3;bcd0<=8; end
			3839: begin bcd3<=3;bcd2<=8;bcd1<=3;bcd0<=9; end
			3840: begin bcd3<=3;bcd2<=8;bcd1<=4;bcd0<=0; end
			3841: begin bcd3<=3;bcd2<=8;bcd1<=4;bcd0<=1; end
			3842: begin bcd3<=3;bcd2<=8;bcd1<=4;bcd0<=2; end
			3843: begin bcd3<=3;bcd2<=8;bcd1<=4;bcd0<=3; end
			3844: begin bcd3<=3;bcd2<=8;bcd1<=4;bcd0<=4; end
			3845: begin bcd3<=3;bcd2<=8;bcd1<=4;bcd0<=5; end
			3846: begin bcd3<=3;bcd2<=8;bcd1<=4;bcd0<=6; end
			3847: begin bcd3<=3;bcd2<=8;bcd1<=4;bcd0<=7; end
			3848: begin bcd3<=3;bcd2<=8;bcd1<=4;bcd0<=8; end
			3849: begin bcd3<=3;bcd2<=8;bcd1<=4;bcd0<=9; end
			3850: begin bcd3<=3;bcd2<=8;bcd1<=5;bcd0<=0; end
			3851: begin bcd3<=3;bcd2<=8;bcd1<=5;bcd0<=1; end
			3852: begin bcd3<=3;bcd2<=8;bcd1<=5;bcd0<=2; end
			3853: begin bcd3<=3;bcd2<=8;bcd1<=5;bcd0<=3; end
			3854: begin bcd3<=3;bcd2<=8;bcd1<=5;bcd0<=4; end
			3855: begin bcd3<=3;bcd2<=8;bcd1<=5;bcd0<=5; end
			3856: begin bcd3<=3;bcd2<=8;bcd1<=5;bcd0<=6; end
			3857: begin bcd3<=3;bcd2<=8;bcd1<=5;bcd0<=7; end
			3858: begin bcd3<=3;bcd2<=8;bcd1<=5;bcd0<=8; end
			3859: begin bcd3<=3;bcd2<=8;bcd1<=5;bcd0<=9; end
			3860: begin bcd3<=3;bcd2<=8;bcd1<=6;bcd0<=0; end
			3861: begin bcd3<=3;bcd2<=8;bcd1<=6;bcd0<=1; end
			3862: begin bcd3<=3;bcd2<=8;bcd1<=6;bcd0<=2; end
			3863: begin bcd3<=3;bcd2<=8;bcd1<=6;bcd0<=3; end
			3864: begin bcd3<=3;bcd2<=8;bcd1<=6;bcd0<=4; end
			3865: begin bcd3<=3;bcd2<=8;bcd1<=6;bcd0<=5; end
			3866: begin bcd3<=3;bcd2<=8;bcd1<=6;bcd0<=6; end
			3867: begin bcd3<=3;bcd2<=8;bcd1<=6;bcd0<=7; end
			3868: begin bcd3<=3;bcd2<=8;bcd1<=6;bcd0<=8; end
			3869: begin bcd3<=3;bcd2<=8;bcd1<=6;bcd0<=9; end
			3870: begin bcd3<=3;bcd2<=8;bcd1<=7;bcd0<=0; end
			3871: begin bcd3<=3;bcd2<=8;bcd1<=7;bcd0<=1; end
			3872: begin bcd3<=3;bcd2<=8;bcd1<=7;bcd0<=2; end
			3873: begin bcd3<=3;bcd2<=8;bcd1<=7;bcd0<=3; end
			3874: begin bcd3<=3;bcd2<=8;bcd1<=7;bcd0<=4; end
			3875: begin bcd3<=3;bcd2<=8;bcd1<=7;bcd0<=5; end
			3876: begin bcd3<=3;bcd2<=8;bcd1<=7;bcd0<=6; end
			3877: begin bcd3<=3;bcd2<=8;bcd1<=7;bcd0<=7; end
			3878: begin bcd3<=3;bcd2<=8;bcd1<=7;bcd0<=8; end
			3879: begin bcd3<=3;bcd2<=8;bcd1<=7;bcd0<=9; end
			3880: begin bcd3<=3;bcd2<=8;bcd1<=8;bcd0<=0; end
			3881: begin bcd3<=3;bcd2<=8;bcd1<=8;bcd0<=1; end
			3882: begin bcd3<=3;bcd2<=8;bcd1<=8;bcd0<=2; end
			3883: begin bcd3<=3;bcd2<=8;bcd1<=8;bcd0<=3; end
			3884: begin bcd3<=3;bcd2<=8;bcd1<=8;bcd0<=4; end
			3885: begin bcd3<=3;bcd2<=8;bcd1<=8;bcd0<=5; end
			3886: begin bcd3<=3;bcd2<=8;bcd1<=8;bcd0<=6; end
			3887: begin bcd3<=3;bcd2<=8;bcd1<=8;bcd0<=7; end
			3888: begin bcd3<=3;bcd2<=8;bcd1<=8;bcd0<=8; end
			3889: begin bcd3<=3;bcd2<=8;bcd1<=8;bcd0<=9; end
			3890: begin bcd3<=3;bcd2<=8;bcd1<=9;bcd0<=0; end
			3891: begin bcd3<=3;bcd2<=8;bcd1<=9;bcd0<=1; end
			3892: begin bcd3<=3;bcd2<=8;bcd1<=9;bcd0<=2; end
			3893: begin bcd3<=3;bcd2<=8;bcd1<=9;bcd0<=3; end
			3894: begin bcd3<=3;bcd2<=8;bcd1<=9;bcd0<=4; end
			3895: begin bcd3<=3;bcd2<=8;bcd1<=9;bcd0<=5; end
			3896: begin bcd3<=3;bcd2<=8;bcd1<=9;bcd0<=6; end
			3897: begin bcd3<=3;bcd2<=8;bcd1<=9;bcd0<=7; end
			3898: begin bcd3<=3;bcd2<=8;bcd1<=9;bcd0<=8; end
			3899: begin bcd3<=3;bcd2<=8;bcd1<=9;bcd0<=9; end
			3900: begin bcd3<=3;bcd2<=9;bcd1<=0;bcd0<=0; end
			3901: begin bcd3<=3;bcd2<=9;bcd1<=0;bcd0<=1; end
			3902: begin bcd3<=3;bcd2<=9;bcd1<=0;bcd0<=2; end
			3903: begin bcd3<=3;bcd2<=9;bcd1<=0;bcd0<=3; end
			3904: begin bcd3<=3;bcd2<=9;bcd1<=0;bcd0<=4; end
			3905: begin bcd3<=3;bcd2<=9;bcd1<=0;bcd0<=5; end
			3906: begin bcd3<=3;bcd2<=9;bcd1<=0;bcd0<=6; end
			3907: begin bcd3<=3;bcd2<=9;bcd1<=0;bcd0<=7; end
			3908: begin bcd3<=3;bcd2<=9;bcd1<=0;bcd0<=8; end
			3909: begin bcd3<=3;bcd2<=9;bcd1<=0;bcd0<=9; end
			3910: begin bcd3<=3;bcd2<=9;bcd1<=1;bcd0<=0; end
			3911: begin bcd3<=3;bcd2<=9;bcd1<=1;bcd0<=1; end
			3912: begin bcd3<=3;bcd2<=9;bcd1<=1;bcd0<=2; end
			3913: begin bcd3<=3;bcd2<=9;bcd1<=1;bcd0<=3; end
			3914: begin bcd3<=3;bcd2<=9;bcd1<=1;bcd0<=4; end
			3915: begin bcd3<=3;bcd2<=9;bcd1<=1;bcd0<=5; end
			3916: begin bcd3<=3;bcd2<=9;bcd1<=1;bcd0<=6; end
			3917: begin bcd3<=3;bcd2<=9;bcd1<=1;bcd0<=7; end
			3918: begin bcd3<=3;bcd2<=9;bcd1<=1;bcd0<=8; end
			3919: begin bcd3<=3;bcd2<=9;bcd1<=1;bcd0<=9; end
			3920: begin bcd3<=3;bcd2<=9;bcd1<=2;bcd0<=0; end
			3921: begin bcd3<=3;bcd2<=9;bcd1<=2;bcd0<=1; end
			3922: begin bcd3<=3;bcd2<=9;bcd1<=2;bcd0<=2; end
			3923: begin bcd3<=3;bcd2<=9;bcd1<=2;bcd0<=3; end
			3924: begin bcd3<=3;bcd2<=9;bcd1<=2;bcd0<=4; end
			3925: begin bcd3<=3;bcd2<=9;bcd1<=2;bcd0<=5; end
			3926: begin bcd3<=3;bcd2<=9;bcd1<=2;bcd0<=6; end
			3927: begin bcd3<=3;bcd2<=9;bcd1<=2;bcd0<=7; end
			3928: begin bcd3<=3;bcd2<=9;bcd1<=2;bcd0<=8; end
			3929: begin bcd3<=3;bcd2<=9;bcd1<=2;bcd0<=9; end
			3930: begin bcd3<=3;bcd2<=9;bcd1<=3;bcd0<=0; end
			3931: begin bcd3<=3;bcd2<=9;bcd1<=3;bcd0<=1; end
			3932: begin bcd3<=3;bcd2<=9;bcd1<=3;bcd0<=2; end
			3933: begin bcd3<=3;bcd2<=9;bcd1<=3;bcd0<=3; end
			3934: begin bcd3<=3;bcd2<=9;bcd1<=3;bcd0<=4; end
			3935: begin bcd3<=3;bcd2<=9;bcd1<=3;bcd0<=5; end
			3936: begin bcd3<=3;bcd2<=9;bcd1<=3;bcd0<=6; end
			3937: begin bcd3<=3;bcd2<=9;bcd1<=3;bcd0<=7; end
			3938: begin bcd3<=3;bcd2<=9;bcd1<=3;bcd0<=8; end
			3939: begin bcd3<=3;bcd2<=9;bcd1<=3;bcd0<=9; end
			3940: begin bcd3<=3;bcd2<=9;bcd1<=4;bcd0<=0; end
			3941: begin bcd3<=3;bcd2<=9;bcd1<=4;bcd0<=1; end
			3942: begin bcd3<=3;bcd2<=9;bcd1<=4;bcd0<=2; end
			3943: begin bcd3<=3;bcd2<=9;bcd1<=4;bcd0<=3; end
			3944: begin bcd3<=3;bcd2<=9;bcd1<=4;bcd0<=4; end
			3945: begin bcd3<=3;bcd2<=9;bcd1<=4;bcd0<=5; end
			3946: begin bcd3<=3;bcd2<=9;bcd1<=4;bcd0<=6; end
			3947: begin bcd3<=3;bcd2<=9;bcd1<=4;bcd0<=7; end
			3948: begin bcd3<=3;bcd2<=9;bcd1<=4;bcd0<=8; end
			3949: begin bcd3<=3;bcd2<=9;bcd1<=4;bcd0<=9; end
			3950: begin bcd3<=3;bcd2<=9;bcd1<=5;bcd0<=0; end
			3951: begin bcd3<=3;bcd2<=9;bcd1<=5;bcd0<=1; end
			3952: begin bcd3<=3;bcd2<=9;bcd1<=5;bcd0<=2; end
			3953: begin bcd3<=3;bcd2<=9;bcd1<=5;bcd0<=3; end
			3954: begin bcd3<=3;bcd2<=9;bcd1<=5;bcd0<=4; end
			3955: begin bcd3<=3;bcd2<=9;bcd1<=5;bcd0<=5; end
			3956: begin bcd3<=3;bcd2<=9;bcd1<=5;bcd0<=6; end
			3957: begin bcd3<=3;bcd2<=9;bcd1<=5;bcd0<=7; end
			3958: begin bcd3<=3;bcd2<=9;bcd1<=5;bcd0<=8; end
			3959: begin bcd3<=3;bcd2<=9;bcd1<=5;bcd0<=9; end
			3960: begin bcd3<=3;bcd2<=9;bcd1<=6;bcd0<=0; end
			3961: begin bcd3<=3;bcd2<=9;bcd1<=6;bcd0<=1; end
			3962: begin bcd3<=3;bcd2<=9;bcd1<=6;bcd0<=2; end
			3963: begin bcd3<=3;bcd2<=9;bcd1<=6;bcd0<=3; end
			3964: begin bcd3<=3;bcd2<=9;bcd1<=6;bcd0<=4; end
			3965: begin bcd3<=3;bcd2<=9;bcd1<=6;bcd0<=5; end
			3966: begin bcd3<=3;bcd2<=9;bcd1<=6;bcd0<=6; end
			3967: begin bcd3<=3;bcd2<=9;bcd1<=6;bcd0<=7; end
			3968: begin bcd3<=3;bcd2<=9;bcd1<=6;bcd0<=8; end
			3969: begin bcd3<=3;bcd2<=9;bcd1<=6;bcd0<=9; end
			3970: begin bcd3<=3;bcd2<=9;bcd1<=7;bcd0<=0; end
			3971: begin bcd3<=3;bcd2<=9;bcd1<=7;bcd0<=1; end
			3972: begin bcd3<=3;bcd2<=9;bcd1<=7;bcd0<=2; end
			3973: begin bcd3<=3;bcd2<=9;bcd1<=7;bcd0<=3; end
			3974: begin bcd3<=3;bcd2<=9;bcd1<=7;bcd0<=4; end
			3975: begin bcd3<=3;bcd2<=9;bcd1<=7;bcd0<=5; end
			3976: begin bcd3<=3;bcd2<=9;bcd1<=7;bcd0<=6; end
			3977: begin bcd3<=3;bcd2<=9;bcd1<=7;bcd0<=7; end
			3978: begin bcd3<=3;bcd2<=9;bcd1<=7;bcd0<=8; end
			3979: begin bcd3<=3;bcd2<=9;bcd1<=7;bcd0<=9; end
			3980: begin bcd3<=3;bcd2<=9;bcd1<=8;bcd0<=0; end
			3981: begin bcd3<=3;bcd2<=9;bcd1<=8;bcd0<=1; end
			3982: begin bcd3<=3;bcd2<=9;bcd1<=8;bcd0<=2; end
			3983: begin bcd3<=3;bcd2<=9;bcd1<=8;bcd0<=3; end
			3984: begin bcd3<=3;bcd2<=9;bcd1<=8;bcd0<=4; end
			3985: begin bcd3<=3;bcd2<=9;bcd1<=8;bcd0<=5; end
			3986: begin bcd3<=3;bcd2<=9;bcd1<=8;bcd0<=6; end
			3987: begin bcd3<=3;bcd2<=9;bcd1<=8;bcd0<=7; end
			3988: begin bcd3<=3;bcd2<=9;bcd1<=8;bcd0<=8; end
			3989: begin bcd3<=3;bcd2<=9;bcd1<=8;bcd0<=9; end
			3990: begin bcd3<=3;bcd2<=9;bcd1<=9;bcd0<=0; end
			3991: begin bcd3<=3;bcd2<=9;bcd1<=9;bcd0<=1; end
			3992: begin bcd3<=3;bcd2<=9;bcd1<=9;bcd0<=2; end
			3993: begin bcd3<=3;bcd2<=9;bcd1<=9;bcd0<=3; end
			3994: begin bcd3<=3;bcd2<=9;bcd1<=9;bcd0<=4; end
			3995: begin bcd3<=3;bcd2<=9;bcd1<=9;bcd0<=5; end
			3996: begin bcd3<=3;bcd2<=9;bcd1<=9;bcd0<=6; end
			3997: begin bcd3<=3;bcd2<=9;bcd1<=9;bcd0<=7; end
			3998: begin bcd3<=3;bcd2<=9;bcd1<=9;bcd0<=8; end
			3999: begin bcd3<=3;bcd2<=9;bcd1<=9;bcd0<=9; end
			4000: begin bcd3<=4;bcd2<=0;bcd1<=0;bcd0<=0; end
			4001: begin bcd3<=4;bcd2<=0;bcd1<=0;bcd0<=1; end
			4002: begin bcd3<=4;bcd2<=0;bcd1<=0;bcd0<=2; end
			4003: begin bcd3<=4;bcd2<=0;bcd1<=0;bcd0<=3; end
			4004: begin bcd3<=4;bcd2<=0;bcd1<=0;bcd0<=4; end
			4005: begin bcd3<=4;bcd2<=0;bcd1<=0;bcd0<=5; end
			4006: begin bcd3<=4;bcd2<=0;bcd1<=0;bcd0<=6; end
			4007: begin bcd3<=4;bcd2<=0;bcd1<=0;bcd0<=7; end
			4008: begin bcd3<=4;bcd2<=0;bcd1<=0;bcd0<=8; end
			4009: begin bcd3<=4;bcd2<=0;bcd1<=0;bcd0<=9; end
			4010: begin bcd3<=4;bcd2<=0;bcd1<=1;bcd0<=0; end
			4011: begin bcd3<=4;bcd2<=0;bcd1<=1;bcd0<=1; end
			4012: begin bcd3<=4;bcd2<=0;bcd1<=1;bcd0<=2; end
			4013: begin bcd3<=4;bcd2<=0;bcd1<=1;bcd0<=3; end
			4014: begin bcd3<=4;bcd2<=0;bcd1<=1;bcd0<=4; end
			4015: begin bcd3<=4;bcd2<=0;bcd1<=1;bcd0<=5; end
			4016: begin bcd3<=4;bcd2<=0;bcd1<=1;bcd0<=6; end
			4017: begin bcd3<=4;bcd2<=0;bcd1<=1;bcd0<=7; end
			4018: begin bcd3<=4;bcd2<=0;bcd1<=1;bcd0<=8; end
			4019: begin bcd3<=4;bcd2<=0;bcd1<=1;bcd0<=9; end
			4020: begin bcd3<=4;bcd2<=0;bcd1<=2;bcd0<=0; end
			4021: begin bcd3<=4;bcd2<=0;bcd1<=2;bcd0<=1; end
			4022: begin bcd3<=4;bcd2<=0;bcd1<=2;bcd0<=2; end
			4023: begin bcd3<=4;bcd2<=0;bcd1<=2;bcd0<=3; end
			4024: begin bcd3<=4;bcd2<=0;bcd1<=2;bcd0<=4; end
			4025: begin bcd3<=4;bcd2<=0;bcd1<=2;bcd0<=5; end
			4026: begin bcd3<=4;bcd2<=0;bcd1<=2;bcd0<=6; end
			4027: begin bcd3<=4;bcd2<=0;bcd1<=2;bcd0<=7; end
			4028: begin bcd3<=4;bcd2<=0;bcd1<=2;bcd0<=8; end
			4029: begin bcd3<=4;bcd2<=0;bcd1<=2;bcd0<=9; end
			4030: begin bcd3<=4;bcd2<=0;bcd1<=3;bcd0<=0; end
			4031: begin bcd3<=4;bcd2<=0;bcd1<=3;bcd0<=1; end
			4032: begin bcd3<=4;bcd2<=0;bcd1<=3;bcd0<=2; end
			4033: begin bcd3<=4;bcd2<=0;bcd1<=3;bcd0<=3; end
			4034: begin bcd3<=4;bcd2<=0;bcd1<=3;bcd0<=4; end
			4035: begin bcd3<=4;bcd2<=0;bcd1<=3;bcd0<=5; end
			4036: begin bcd3<=4;bcd2<=0;bcd1<=3;bcd0<=6; end
			4037: begin bcd3<=4;bcd2<=0;bcd1<=3;bcd0<=7; end
			4038: begin bcd3<=4;bcd2<=0;bcd1<=3;bcd0<=8; end
			4039: begin bcd3<=4;bcd2<=0;bcd1<=3;bcd0<=9; end
			4040: begin bcd3<=4;bcd2<=0;bcd1<=4;bcd0<=0; end
			4041: begin bcd3<=4;bcd2<=0;bcd1<=4;bcd0<=1; end
			4042: begin bcd3<=4;bcd2<=0;bcd1<=4;bcd0<=2; end
			4043: begin bcd3<=4;bcd2<=0;bcd1<=4;bcd0<=3; end
			4044: begin bcd3<=4;bcd2<=0;bcd1<=4;bcd0<=4; end
			4045: begin bcd3<=4;bcd2<=0;bcd1<=4;bcd0<=5; end
			4046: begin bcd3<=4;bcd2<=0;bcd1<=4;bcd0<=6; end
			4047: begin bcd3<=4;bcd2<=0;bcd1<=4;bcd0<=7; end
			4048: begin bcd3<=4;bcd2<=0;bcd1<=4;bcd0<=8; end
			4049: begin bcd3<=4;bcd2<=0;bcd1<=4;bcd0<=9; end
			4050: begin bcd3<=4;bcd2<=0;bcd1<=5;bcd0<=0; end
			4051: begin bcd3<=4;bcd2<=0;bcd1<=5;bcd0<=1; end
			4052: begin bcd3<=4;bcd2<=0;bcd1<=5;bcd0<=2; end
			4053: begin bcd3<=4;bcd2<=0;bcd1<=5;bcd0<=3; end
			4054: begin bcd3<=4;bcd2<=0;bcd1<=5;bcd0<=4; end
			4055: begin bcd3<=4;bcd2<=0;bcd1<=5;bcd0<=5; end
			4056: begin bcd3<=4;bcd2<=0;bcd1<=5;bcd0<=6; end
			4057: begin bcd3<=4;bcd2<=0;bcd1<=5;bcd0<=7; end
			4058: begin bcd3<=4;bcd2<=0;bcd1<=5;bcd0<=8; end
			4059: begin bcd3<=4;bcd2<=0;bcd1<=5;bcd0<=9; end
			4060: begin bcd3<=4;bcd2<=0;bcd1<=6;bcd0<=0; end
			4061: begin bcd3<=4;bcd2<=0;bcd1<=6;bcd0<=1; end
			4062: begin bcd3<=4;bcd2<=0;bcd1<=6;bcd0<=2; end
			4063: begin bcd3<=4;bcd2<=0;bcd1<=6;bcd0<=3; end
			4064: begin bcd3<=4;bcd2<=0;bcd1<=6;bcd0<=4; end
			4065: begin bcd3<=4;bcd2<=0;bcd1<=6;bcd0<=5; end
			4066: begin bcd3<=4;bcd2<=0;bcd1<=6;bcd0<=6; end
			4067: begin bcd3<=4;bcd2<=0;bcd1<=6;bcd0<=7; end
			4068: begin bcd3<=4;bcd2<=0;bcd1<=6;bcd0<=8; end
			4069: begin bcd3<=4;bcd2<=0;bcd1<=6;bcd0<=9; end
			4070: begin bcd3<=4;bcd2<=0;bcd1<=7;bcd0<=0; end
			4071: begin bcd3<=4;bcd2<=0;bcd1<=7;bcd0<=1; end
			4072: begin bcd3<=4;bcd2<=0;bcd1<=7;bcd0<=2; end
			4073: begin bcd3<=4;bcd2<=0;bcd1<=7;bcd0<=3; end
			4074: begin bcd3<=4;bcd2<=0;bcd1<=7;bcd0<=4; end
			4075: begin bcd3<=4;bcd2<=0;bcd1<=7;bcd0<=5; end
			4076: begin bcd3<=4;bcd2<=0;bcd1<=7;bcd0<=6; end
			4077: begin bcd3<=4;bcd2<=0;bcd1<=7;bcd0<=7; end
			4078: begin bcd3<=4;bcd2<=0;bcd1<=7;bcd0<=8; end
			4079: begin bcd3<=4;bcd2<=0;bcd1<=7;bcd0<=9; end
			4080: begin bcd3<=4;bcd2<=0;bcd1<=8;bcd0<=0; end
			4081: begin bcd3<=4;bcd2<=0;bcd1<=8;bcd0<=1; end
			4082: begin bcd3<=4;bcd2<=0;bcd1<=8;bcd0<=2; end
			4083: begin bcd3<=4;bcd2<=0;bcd1<=8;bcd0<=3; end
			4084: begin bcd3<=4;bcd2<=0;bcd1<=8;bcd0<=4; end
			4085: begin bcd3<=4;bcd2<=0;bcd1<=8;bcd0<=5; end
			4086: begin bcd3<=4;bcd2<=0;bcd1<=8;bcd0<=6; end
			4087: begin bcd3<=4;bcd2<=0;bcd1<=8;bcd0<=7; end
			4088: begin bcd3<=4;bcd2<=0;bcd1<=8;bcd0<=8; end
			4089: begin bcd3<=4;bcd2<=0;bcd1<=8;bcd0<=9; end
			4090: begin bcd3<=4;bcd2<=0;bcd1<=9;bcd0<=0; end
			4091: begin bcd3<=4;bcd2<=0;bcd1<=9;bcd0<=1; end
			4092: begin bcd3<=4;bcd2<=0;bcd1<=9;bcd0<=2; end
			4093: begin bcd3<=4;bcd2<=0;bcd1<=9;bcd0<=3; end
			4094: begin bcd3<=4;bcd2<=0;bcd1<=9;bcd0<=4; end
			4095: begin bcd3<=4;bcd2<=0;bcd1<=9;bcd0<=5; end
			4096: begin bcd3<=4;bcd2<=0;bcd1<=9;bcd0<=6; end
			4097: begin bcd3<=4;bcd2<=0;bcd1<=9;bcd0<=7; end
			4098: begin bcd3<=4;bcd2<=0;bcd1<=9;bcd0<=8; end
			4099: begin bcd3<=4;bcd2<=0;bcd1<=9;bcd0<=9; end
			4100: begin bcd3<=4;bcd2<=1;bcd1<=0;bcd0<=0; end
			4101: begin bcd3<=4;bcd2<=1;bcd1<=0;bcd0<=1; end
			4102: begin bcd3<=4;bcd2<=1;bcd1<=0;bcd0<=2; end
			4103: begin bcd3<=4;bcd2<=1;bcd1<=0;bcd0<=3; end
			4104: begin bcd3<=4;bcd2<=1;bcd1<=0;bcd0<=4; end
			4105: begin bcd3<=4;bcd2<=1;bcd1<=0;bcd0<=5; end
			4106: begin bcd3<=4;bcd2<=1;bcd1<=0;bcd0<=6; end
			4107: begin bcd3<=4;bcd2<=1;bcd1<=0;bcd0<=7; end
			4108: begin bcd3<=4;bcd2<=1;bcd1<=0;bcd0<=8; end
			4109: begin bcd3<=4;bcd2<=1;bcd1<=0;bcd0<=9; end
			4110: begin bcd3<=4;bcd2<=1;bcd1<=1;bcd0<=0; end
			4111: begin bcd3<=4;bcd2<=1;bcd1<=1;bcd0<=1; end
			4112: begin bcd3<=4;bcd2<=1;bcd1<=1;bcd0<=2; end
			4113: begin bcd3<=4;bcd2<=1;bcd1<=1;bcd0<=3; end
			4114: begin bcd3<=4;bcd2<=1;bcd1<=1;bcd0<=4; end
			4115: begin bcd3<=4;bcd2<=1;bcd1<=1;bcd0<=5; end
			4116: begin bcd3<=4;bcd2<=1;bcd1<=1;bcd0<=6; end
			4117: begin bcd3<=4;bcd2<=1;bcd1<=1;bcd0<=7; end
			4118: begin bcd3<=4;bcd2<=1;bcd1<=1;bcd0<=8; end
			4119: begin bcd3<=4;bcd2<=1;bcd1<=1;bcd0<=9; end
			4120: begin bcd3<=4;bcd2<=1;bcd1<=2;bcd0<=0; end
			4121: begin bcd3<=4;bcd2<=1;bcd1<=2;bcd0<=1; end
			4122: begin bcd3<=4;bcd2<=1;bcd1<=2;bcd0<=2; end
			4123: begin bcd3<=4;bcd2<=1;bcd1<=2;bcd0<=3; end
			4124: begin bcd3<=4;bcd2<=1;bcd1<=2;bcd0<=4; end
			4125: begin bcd3<=4;bcd2<=1;bcd1<=2;bcd0<=5; end
			4126: begin bcd3<=4;bcd2<=1;bcd1<=2;bcd0<=6; end
			4127: begin bcd3<=4;bcd2<=1;bcd1<=2;bcd0<=7; end
			4128: begin bcd3<=4;bcd2<=1;bcd1<=2;bcd0<=8; end
			4129: begin bcd3<=4;bcd2<=1;bcd1<=2;bcd0<=9; end
			4130: begin bcd3<=4;bcd2<=1;bcd1<=3;bcd0<=0; end
			4131: begin bcd3<=4;bcd2<=1;bcd1<=3;bcd0<=1; end
			4132: begin bcd3<=4;bcd2<=1;bcd1<=3;bcd0<=2; end
			4133: begin bcd3<=4;bcd2<=1;bcd1<=3;bcd0<=3; end
			4134: begin bcd3<=4;bcd2<=1;bcd1<=3;bcd0<=4; end
			4135: begin bcd3<=4;bcd2<=1;bcd1<=3;bcd0<=5; end
			4136: begin bcd3<=4;bcd2<=1;bcd1<=3;bcd0<=6; end
			4137: begin bcd3<=4;bcd2<=1;bcd1<=3;bcd0<=7; end
			4138: begin bcd3<=4;bcd2<=1;bcd1<=3;bcd0<=8; end
			4139: begin bcd3<=4;bcd2<=1;bcd1<=3;bcd0<=9; end
			4140: begin bcd3<=4;bcd2<=1;bcd1<=4;bcd0<=0; end
			4141: begin bcd3<=4;bcd2<=1;bcd1<=4;bcd0<=1; end
			4142: begin bcd3<=4;bcd2<=1;bcd1<=4;bcd0<=2; end
			4143: begin bcd3<=4;bcd2<=1;bcd1<=4;bcd0<=3; end
			4144: begin bcd3<=4;bcd2<=1;bcd1<=4;bcd0<=4; end
			4145: begin bcd3<=4;bcd2<=1;bcd1<=4;bcd0<=5; end
			4146: begin bcd3<=4;bcd2<=1;bcd1<=4;bcd0<=6; end
			4147: begin bcd3<=4;bcd2<=1;bcd1<=4;bcd0<=7; end
			4148: begin bcd3<=4;bcd2<=1;bcd1<=4;bcd0<=8; end
			4149: begin bcd3<=4;bcd2<=1;bcd1<=4;bcd0<=9; end
			4150: begin bcd3<=4;bcd2<=1;bcd1<=5;bcd0<=0; end
			4151: begin bcd3<=4;bcd2<=1;bcd1<=5;bcd0<=1; end
			4152: begin bcd3<=4;bcd2<=1;bcd1<=5;bcd0<=2; end
			4153: begin bcd3<=4;bcd2<=1;bcd1<=5;bcd0<=3; end
			4154: begin bcd3<=4;bcd2<=1;bcd1<=5;bcd0<=4; end
			4155: begin bcd3<=4;bcd2<=1;bcd1<=5;bcd0<=5; end
			4156: begin bcd3<=4;bcd2<=1;bcd1<=5;bcd0<=6; end
			4157: begin bcd3<=4;bcd2<=1;bcd1<=5;bcd0<=7; end
			4158: begin bcd3<=4;bcd2<=1;bcd1<=5;bcd0<=8; end
			4159: begin bcd3<=4;bcd2<=1;bcd1<=5;bcd0<=9; end
			4160: begin bcd3<=4;bcd2<=1;bcd1<=6;bcd0<=0; end
			4161: begin bcd3<=4;bcd2<=1;bcd1<=6;bcd0<=1; end
			4162: begin bcd3<=4;bcd2<=1;bcd1<=6;bcd0<=2; end
			4163: begin bcd3<=4;bcd2<=1;bcd1<=6;bcd0<=3; end
			4164: begin bcd3<=4;bcd2<=1;bcd1<=6;bcd0<=4; end
			4165: begin bcd3<=4;bcd2<=1;bcd1<=6;bcd0<=5; end
			4166: begin bcd3<=4;bcd2<=1;bcd1<=6;bcd0<=6; end
			4167: begin bcd3<=4;bcd2<=1;bcd1<=6;bcd0<=7; end
			4168: begin bcd3<=4;bcd2<=1;bcd1<=6;bcd0<=8; end
			4169: begin bcd3<=4;bcd2<=1;bcd1<=6;bcd0<=9; end
			4170: begin bcd3<=4;bcd2<=1;bcd1<=7;bcd0<=0; end
			4171: begin bcd3<=4;bcd2<=1;bcd1<=7;bcd0<=1; end
			4172: begin bcd3<=4;bcd2<=1;bcd1<=7;bcd0<=2; end
			4173: begin bcd3<=4;bcd2<=1;bcd1<=7;bcd0<=3; end
			4174: begin bcd3<=4;bcd2<=1;bcd1<=7;bcd0<=4; end
			4175: begin bcd3<=4;bcd2<=1;bcd1<=7;bcd0<=5; end
			4176: begin bcd3<=4;bcd2<=1;bcd1<=7;bcd0<=6; end
			4177: begin bcd3<=4;bcd2<=1;bcd1<=7;bcd0<=7; end
			4178: begin bcd3<=4;bcd2<=1;bcd1<=7;bcd0<=8; end
			4179: begin bcd3<=4;bcd2<=1;bcd1<=7;bcd0<=9; end
			4180: begin bcd3<=4;bcd2<=1;bcd1<=8;bcd0<=0; end
			4181: begin bcd3<=4;bcd2<=1;bcd1<=8;bcd0<=1; end
			4182: begin bcd3<=4;bcd2<=1;bcd1<=8;bcd0<=2; end
			4183: begin bcd3<=4;bcd2<=1;bcd1<=8;bcd0<=3; end
			4184: begin bcd3<=4;bcd2<=1;bcd1<=8;bcd0<=4; end
			4185: begin bcd3<=4;bcd2<=1;bcd1<=8;bcd0<=5; end
			4186: begin bcd3<=4;bcd2<=1;bcd1<=8;bcd0<=6; end
			4187: begin bcd3<=4;bcd2<=1;bcd1<=8;bcd0<=7; end
			4188: begin bcd3<=4;bcd2<=1;bcd1<=8;bcd0<=8; end
			4189: begin bcd3<=4;bcd2<=1;bcd1<=8;bcd0<=9; end
			4190: begin bcd3<=4;bcd2<=1;bcd1<=9;bcd0<=0; end
			4191: begin bcd3<=4;bcd2<=1;bcd1<=9;bcd0<=1; end
			4192: begin bcd3<=4;bcd2<=1;bcd1<=9;bcd0<=2; end
			4193: begin bcd3<=4;bcd2<=1;bcd1<=9;bcd0<=3; end
			4194: begin bcd3<=4;bcd2<=1;bcd1<=9;bcd0<=4; end
			4195: begin bcd3<=4;bcd2<=1;bcd1<=9;bcd0<=5; end
			4196: begin bcd3<=4;bcd2<=1;bcd1<=9;bcd0<=6; end
			4197: begin bcd3<=4;bcd2<=1;bcd1<=9;bcd0<=7; end
			4198: begin bcd3<=4;bcd2<=1;bcd1<=9;bcd0<=8; end
			4199: begin bcd3<=4;bcd2<=1;bcd1<=9;bcd0<=9; end
			4200: begin bcd3<=4;bcd2<=2;bcd1<=0;bcd0<=0; end
			4201: begin bcd3<=4;bcd2<=2;bcd1<=0;bcd0<=1; end
			4202: begin bcd3<=4;bcd2<=2;bcd1<=0;bcd0<=2; end
			4203: begin bcd3<=4;bcd2<=2;bcd1<=0;bcd0<=3; end
			4204: begin bcd3<=4;bcd2<=2;bcd1<=0;bcd0<=4; end
			4205: begin bcd3<=4;bcd2<=2;bcd1<=0;bcd0<=5; end
			4206: begin bcd3<=4;bcd2<=2;bcd1<=0;bcd0<=6; end
			4207: begin bcd3<=4;bcd2<=2;bcd1<=0;bcd0<=7; end
			4208: begin bcd3<=4;bcd2<=2;bcd1<=0;bcd0<=8; end
			4209: begin bcd3<=4;bcd2<=2;bcd1<=0;bcd0<=9; end
			4210: begin bcd3<=4;bcd2<=2;bcd1<=1;bcd0<=0; end
			4211: begin bcd3<=4;bcd2<=2;bcd1<=1;bcd0<=1; end
			4212: begin bcd3<=4;bcd2<=2;bcd1<=1;bcd0<=2; end
			4213: begin bcd3<=4;bcd2<=2;bcd1<=1;bcd0<=3; end
			4214: begin bcd3<=4;bcd2<=2;bcd1<=1;bcd0<=4; end
			4215: begin bcd3<=4;bcd2<=2;bcd1<=1;bcd0<=5; end
			4216: begin bcd3<=4;bcd2<=2;bcd1<=1;bcd0<=6; end
			4217: begin bcd3<=4;bcd2<=2;bcd1<=1;bcd0<=7; end
			4218: begin bcd3<=4;bcd2<=2;bcd1<=1;bcd0<=8; end
			4219: begin bcd3<=4;bcd2<=2;bcd1<=1;bcd0<=9; end
			4220: begin bcd3<=4;bcd2<=2;bcd1<=2;bcd0<=0; end
			4221: begin bcd3<=4;bcd2<=2;bcd1<=2;bcd0<=1; end
			4222: begin bcd3<=4;bcd2<=2;bcd1<=2;bcd0<=2; end
			4223: begin bcd3<=4;bcd2<=2;bcd1<=2;bcd0<=3; end
			4224: begin bcd3<=4;bcd2<=2;bcd1<=2;bcd0<=4; end
			4225: begin bcd3<=4;bcd2<=2;bcd1<=2;bcd0<=5; end
			4226: begin bcd3<=4;bcd2<=2;bcd1<=2;bcd0<=6; end
			4227: begin bcd3<=4;bcd2<=2;bcd1<=2;bcd0<=7; end
			4228: begin bcd3<=4;bcd2<=2;bcd1<=2;bcd0<=8; end
			4229: begin bcd3<=4;bcd2<=2;bcd1<=2;bcd0<=9; end
			4230: begin bcd3<=4;bcd2<=2;bcd1<=3;bcd0<=0; end
			4231: begin bcd3<=4;bcd2<=2;bcd1<=3;bcd0<=1; end
			4232: begin bcd3<=4;bcd2<=2;bcd1<=3;bcd0<=2; end
			4233: begin bcd3<=4;bcd2<=2;bcd1<=3;bcd0<=3; end
			4234: begin bcd3<=4;bcd2<=2;bcd1<=3;bcd0<=4; end
			4235: begin bcd3<=4;bcd2<=2;bcd1<=3;bcd0<=5; end
			4236: begin bcd3<=4;bcd2<=2;bcd1<=3;bcd0<=6; end
			4237: begin bcd3<=4;bcd2<=2;bcd1<=3;bcd0<=7; end
			4238: begin bcd3<=4;bcd2<=2;bcd1<=3;bcd0<=8; end
			4239: begin bcd3<=4;bcd2<=2;bcd1<=3;bcd0<=9; end
			4240: begin bcd3<=4;bcd2<=2;bcd1<=4;bcd0<=0; end
			4241: begin bcd3<=4;bcd2<=2;bcd1<=4;bcd0<=1; end
			4242: begin bcd3<=4;bcd2<=2;bcd1<=4;bcd0<=2; end
			4243: begin bcd3<=4;bcd2<=2;bcd1<=4;bcd0<=3; end
			4244: begin bcd3<=4;bcd2<=2;bcd1<=4;bcd0<=4; end
			4245: begin bcd3<=4;bcd2<=2;bcd1<=4;bcd0<=5; end
			4246: begin bcd3<=4;bcd2<=2;bcd1<=4;bcd0<=6; end
			4247: begin bcd3<=4;bcd2<=2;bcd1<=4;bcd0<=7; end
			4248: begin bcd3<=4;bcd2<=2;bcd1<=4;bcd0<=8; end
			4249: begin bcd3<=4;bcd2<=2;bcd1<=4;bcd0<=9; end
			4250: begin bcd3<=4;bcd2<=2;bcd1<=5;bcd0<=0; end
			4251: begin bcd3<=4;bcd2<=2;bcd1<=5;bcd0<=1; end
			4252: begin bcd3<=4;bcd2<=2;bcd1<=5;bcd0<=2; end
			4253: begin bcd3<=4;bcd2<=2;bcd1<=5;bcd0<=3; end
			4254: begin bcd3<=4;bcd2<=2;bcd1<=5;bcd0<=4; end
			4255: begin bcd3<=4;bcd2<=2;bcd1<=5;bcd0<=5; end
			4256: begin bcd3<=4;bcd2<=2;bcd1<=5;bcd0<=6; end
			4257: begin bcd3<=4;bcd2<=2;bcd1<=5;bcd0<=7; end
			4258: begin bcd3<=4;bcd2<=2;bcd1<=5;bcd0<=8; end
			4259: begin bcd3<=4;bcd2<=2;bcd1<=5;bcd0<=9; end
			4260: begin bcd3<=4;bcd2<=2;bcd1<=6;bcd0<=0; end
			4261: begin bcd3<=4;bcd2<=2;bcd1<=6;bcd0<=1; end
			4262: begin bcd3<=4;bcd2<=2;bcd1<=6;bcd0<=2; end
			4263: begin bcd3<=4;bcd2<=2;bcd1<=6;bcd0<=3; end
			4264: begin bcd3<=4;bcd2<=2;bcd1<=6;bcd0<=4; end
			4265: begin bcd3<=4;bcd2<=2;bcd1<=6;bcd0<=5; end
			4266: begin bcd3<=4;bcd2<=2;bcd1<=6;bcd0<=6; end
			4267: begin bcd3<=4;bcd2<=2;bcd1<=6;bcd0<=7; end
			4268: begin bcd3<=4;bcd2<=2;bcd1<=6;bcd0<=8; end
			4269: begin bcd3<=4;bcd2<=2;bcd1<=6;bcd0<=9; end
			4270: begin bcd3<=4;bcd2<=2;bcd1<=7;bcd0<=0; end
			4271: begin bcd3<=4;bcd2<=2;bcd1<=7;bcd0<=1; end
			4272: begin bcd3<=4;bcd2<=2;bcd1<=7;bcd0<=2; end
			4273: begin bcd3<=4;bcd2<=2;bcd1<=7;bcd0<=3; end
			4274: begin bcd3<=4;bcd2<=2;bcd1<=7;bcd0<=4; end
			4275: begin bcd3<=4;bcd2<=2;bcd1<=7;bcd0<=5; end
			4276: begin bcd3<=4;bcd2<=2;bcd1<=7;bcd0<=6; end
			4277: begin bcd3<=4;bcd2<=2;bcd1<=7;bcd0<=7; end
			4278: begin bcd3<=4;bcd2<=2;bcd1<=7;bcd0<=8; end
			4279: begin bcd3<=4;bcd2<=2;bcd1<=7;bcd0<=9; end
			4280: begin bcd3<=4;bcd2<=2;bcd1<=8;bcd0<=0; end
			4281: begin bcd3<=4;bcd2<=2;bcd1<=8;bcd0<=1; end
			4282: begin bcd3<=4;bcd2<=2;bcd1<=8;bcd0<=2; end
			4283: begin bcd3<=4;bcd2<=2;bcd1<=8;bcd0<=3; end
			4284: begin bcd3<=4;bcd2<=2;bcd1<=8;bcd0<=4; end
			4285: begin bcd3<=4;bcd2<=2;bcd1<=8;bcd0<=5; end
			4286: begin bcd3<=4;bcd2<=2;bcd1<=8;bcd0<=6; end
			4287: begin bcd3<=4;bcd2<=2;bcd1<=8;bcd0<=7; end
			4288: begin bcd3<=4;bcd2<=2;bcd1<=8;bcd0<=8; end
			4289: begin bcd3<=4;bcd2<=2;bcd1<=8;bcd0<=9; end
			4290: begin bcd3<=4;bcd2<=2;bcd1<=9;bcd0<=0; end
			4291: begin bcd3<=4;bcd2<=2;bcd1<=9;bcd0<=1; end
			4292: begin bcd3<=4;bcd2<=2;bcd1<=9;bcd0<=2; end
			4293: begin bcd3<=4;bcd2<=2;bcd1<=9;bcd0<=3; end
			4294: begin bcd3<=4;bcd2<=2;bcd1<=9;bcd0<=4; end
			4295: begin bcd3<=4;bcd2<=2;bcd1<=9;bcd0<=5; end
			4296: begin bcd3<=4;bcd2<=2;bcd1<=9;bcd0<=6; end
			4297: begin bcd3<=4;bcd2<=2;bcd1<=9;bcd0<=7; end
			4298: begin bcd3<=4;bcd2<=2;bcd1<=9;bcd0<=8; end
			4299: begin bcd3<=4;bcd2<=2;bcd1<=9;bcd0<=9; end
			4300: begin bcd3<=4;bcd2<=3;bcd1<=0;bcd0<=0; end
			4301: begin bcd3<=4;bcd2<=3;bcd1<=0;bcd0<=1; end
			4302: begin bcd3<=4;bcd2<=3;bcd1<=0;bcd0<=2; end
			4303: begin bcd3<=4;bcd2<=3;bcd1<=0;bcd0<=3; end
			4304: begin bcd3<=4;bcd2<=3;bcd1<=0;bcd0<=4; end
			4305: begin bcd3<=4;bcd2<=3;bcd1<=0;bcd0<=5; end
			4306: begin bcd3<=4;bcd2<=3;bcd1<=0;bcd0<=6; end
			4307: begin bcd3<=4;bcd2<=3;bcd1<=0;bcd0<=7; end
			4308: begin bcd3<=4;bcd2<=3;bcd1<=0;bcd0<=8; end
			4309: begin bcd3<=4;bcd2<=3;bcd1<=0;bcd0<=9; end
			4310: begin bcd3<=4;bcd2<=3;bcd1<=1;bcd0<=0; end
			4311: begin bcd3<=4;bcd2<=3;bcd1<=1;bcd0<=1; end
			4312: begin bcd3<=4;bcd2<=3;bcd1<=1;bcd0<=2; end
			4313: begin bcd3<=4;bcd2<=3;bcd1<=1;bcd0<=3; end
			4314: begin bcd3<=4;bcd2<=3;bcd1<=1;bcd0<=4; end
			4315: begin bcd3<=4;bcd2<=3;bcd1<=1;bcd0<=5; end
			4316: begin bcd3<=4;bcd2<=3;bcd1<=1;bcd0<=6; end
			4317: begin bcd3<=4;bcd2<=3;bcd1<=1;bcd0<=7; end
			4318: begin bcd3<=4;bcd2<=3;bcd1<=1;bcd0<=8; end
			4319: begin bcd3<=4;bcd2<=3;bcd1<=1;bcd0<=9; end
			4320: begin bcd3<=4;bcd2<=3;bcd1<=2;bcd0<=0; end
			4321: begin bcd3<=4;bcd2<=3;bcd1<=2;bcd0<=1; end
			4322: begin bcd3<=4;bcd2<=3;bcd1<=2;bcd0<=2; end
			4323: begin bcd3<=4;bcd2<=3;bcd1<=2;bcd0<=3; end
			4324: begin bcd3<=4;bcd2<=3;bcd1<=2;bcd0<=4; end
			4325: begin bcd3<=4;bcd2<=3;bcd1<=2;bcd0<=5; end
			4326: begin bcd3<=4;bcd2<=3;bcd1<=2;bcd0<=6; end
			4327: begin bcd3<=4;bcd2<=3;bcd1<=2;bcd0<=7; end
			4328: begin bcd3<=4;bcd2<=3;bcd1<=2;bcd0<=8; end
			4329: begin bcd3<=4;bcd2<=3;bcd1<=2;bcd0<=9; end
			4330: begin bcd3<=4;bcd2<=3;bcd1<=3;bcd0<=0; end
			4331: begin bcd3<=4;bcd2<=3;bcd1<=3;bcd0<=1; end
			4332: begin bcd3<=4;bcd2<=3;bcd1<=3;bcd0<=2; end
			4333: begin bcd3<=4;bcd2<=3;bcd1<=3;bcd0<=3; end
			4334: begin bcd3<=4;bcd2<=3;bcd1<=3;bcd0<=4; end
			4335: begin bcd3<=4;bcd2<=3;bcd1<=3;bcd0<=5; end
			4336: begin bcd3<=4;bcd2<=3;bcd1<=3;bcd0<=6; end
			4337: begin bcd3<=4;bcd2<=3;bcd1<=3;bcd0<=7; end
			4338: begin bcd3<=4;bcd2<=3;bcd1<=3;bcd0<=8; end
			4339: begin bcd3<=4;bcd2<=3;bcd1<=3;bcd0<=9; end
			4340: begin bcd3<=4;bcd2<=3;bcd1<=4;bcd0<=0; end
			4341: begin bcd3<=4;bcd2<=3;bcd1<=4;bcd0<=1; end
			4342: begin bcd3<=4;bcd2<=3;bcd1<=4;bcd0<=2; end
			4343: begin bcd3<=4;bcd2<=3;bcd1<=4;bcd0<=3; end
			4344: begin bcd3<=4;bcd2<=3;bcd1<=4;bcd0<=4; end
			4345: begin bcd3<=4;bcd2<=3;bcd1<=4;bcd0<=5; end
			4346: begin bcd3<=4;bcd2<=3;bcd1<=4;bcd0<=6; end
			4347: begin bcd3<=4;bcd2<=3;bcd1<=4;bcd0<=7; end
			4348: begin bcd3<=4;bcd2<=3;bcd1<=4;bcd0<=8; end
			4349: begin bcd3<=4;bcd2<=3;bcd1<=4;bcd0<=9; end
			4350: begin bcd3<=4;bcd2<=3;bcd1<=5;bcd0<=0; end
			4351: begin bcd3<=4;bcd2<=3;bcd1<=5;bcd0<=1; end
			4352: begin bcd3<=4;bcd2<=3;bcd1<=5;bcd0<=2; end
			4353: begin bcd3<=4;bcd2<=3;bcd1<=5;bcd0<=3; end
			4354: begin bcd3<=4;bcd2<=3;bcd1<=5;bcd0<=4; end
			4355: begin bcd3<=4;bcd2<=3;bcd1<=5;bcd0<=5; end
			4356: begin bcd3<=4;bcd2<=3;bcd1<=5;bcd0<=6; end
			4357: begin bcd3<=4;bcd2<=3;bcd1<=5;bcd0<=7; end
			4358: begin bcd3<=4;bcd2<=3;bcd1<=5;bcd0<=8; end
			4359: begin bcd3<=4;bcd2<=3;bcd1<=5;bcd0<=9; end
			4360: begin bcd3<=4;bcd2<=3;bcd1<=6;bcd0<=0; end
			4361: begin bcd3<=4;bcd2<=3;bcd1<=6;bcd0<=1; end
			4362: begin bcd3<=4;bcd2<=3;bcd1<=6;bcd0<=2; end
			4363: begin bcd3<=4;bcd2<=3;bcd1<=6;bcd0<=3; end
			4364: begin bcd3<=4;bcd2<=3;bcd1<=6;bcd0<=4; end
			4365: begin bcd3<=4;bcd2<=3;bcd1<=6;bcd0<=5; end
			4366: begin bcd3<=4;bcd2<=3;bcd1<=6;bcd0<=6; end
			4367: begin bcd3<=4;bcd2<=3;bcd1<=6;bcd0<=7; end
			4368: begin bcd3<=4;bcd2<=3;bcd1<=6;bcd0<=8; end
			4369: begin bcd3<=4;bcd2<=3;bcd1<=6;bcd0<=9; end
			4370: begin bcd3<=4;bcd2<=3;bcd1<=7;bcd0<=0; end
			4371: begin bcd3<=4;bcd2<=3;bcd1<=7;bcd0<=1; end
			4372: begin bcd3<=4;bcd2<=3;bcd1<=7;bcd0<=2; end
			4373: begin bcd3<=4;bcd2<=3;bcd1<=7;bcd0<=3; end
			4374: begin bcd3<=4;bcd2<=3;bcd1<=7;bcd0<=4; end
			4375: begin bcd3<=4;bcd2<=3;bcd1<=7;bcd0<=5; end
			4376: begin bcd3<=4;bcd2<=3;bcd1<=7;bcd0<=6; end
			4377: begin bcd3<=4;bcd2<=3;bcd1<=7;bcd0<=7; end
			4378: begin bcd3<=4;bcd2<=3;bcd1<=7;bcd0<=8; end
			4379: begin bcd3<=4;bcd2<=3;bcd1<=7;bcd0<=9; end
			4380: begin bcd3<=4;bcd2<=3;bcd1<=8;bcd0<=0; end
			4381: begin bcd3<=4;bcd2<=3;bcd1<=8;bcd0<=1; end
			4382: begin bcd3<=4;bcd2<=3;bcd1<=8;bcd0<=2; end
			4383: begin bcd3<=4;bcd2<=3;bcd1<=8;bcd0<=3; end
			4384: begin bcd3<=4;bcd2<=3;bcd1<=8;bcd0<=4; end
			4385: begin bcd3<=4;bcd2<=3;bcd1<=8;bcd0<=5; end
			4386: begin bcd3<=4;bcd2<=3;bcd1<=8;bcd0<=6; end
			4387: begin bcd3<=4;bcd2<=3;bcd1<=8;bcd0<=7; end
			4388: begin bcd3<=4;bcd2<=3;bcd1<=8;bcd0<=8; end
			4389: begin bcd3<=4;bcd2<=3;bcd1<=8;bcd0<=9; end
			4390: begin bcd3<=4;bcd2<=3;bcd1<=9;bcd0<=0; end
			4391: begin bcd3<=4;bcd2<=3;bcd1<=9;bcd0<=1; end
			4392: begin bcd3<=4;bcd2<=3;bcd1<=9;bcd0<=2; end
			4393: begin bcd3<=4;bcd2<=3;bcd1<=9;bcd0<=3; end
			4394: begin bcd3<=4;bcd2<=3;bcd1<=9;bcd0<=4; end
			4395: begin bcd3<=4;bcd2<=3;bcd1<=9;bcd0<=5; end
			4396: begin bcd3<=4;bcd2<=3;bcd1<=9;bcd0<=6; end
			4397: begin bcd3<=4;bcd2<=3;bcd1<=9;bcd0<=7; end
			4398: begin bcd3<=4;bcd2<=3;bcd1<=9;bcd0<=8; end
			4399: begin bcd3<=4;bcd2<=3;bcd1<=9;bcd0<=9; end
			4400: begin bcd3<=4;bcd2<=4;bcd1<=0;bcd0<=0; end
			4401: begin bcd3<=4;bcd2<=4;bcd1<=0;bcd0<=1; end
			4402: begin bcd3<=4;bcd2<=4;bcd1<=0;bcd0<=2; end
			4403: begin bcd3<=4;bcd2<=4;bcd1<=0;bcd0<=3; end
			4404: begin bcd3<=4;bcd2<=4;bcd1<=0;bcd0<=4; end
			4405: begin bcd3<=4;bcd2<=4;bcd1<=0;bcd0<=5; end
			4406: begin bcd3<=4;bcd2<=4;bcd1<=0;bcd0<=6; end
			4407: begin bcd3<=4;bcd2<=4;bcd1<=0;bcd0<=7; end
			4408: begin bcd3<=4;bcd2<=4;bcd1<=0;bcd0<=8; end
			4409: begin bcd3<=4;bcd2<=4;bcd1<=0;bcd0<=9; end
			4410: begin bcd3<=4;bcd2<=4;bcd1<=1;bcd0<=0; end
			4411: begin bcd3<=4;bcd2<=4;bcd1<=1;bcd0<=1; end
			4412: begin bcd3<=4;bcd2<=4;bcd1<=1;bcd0<=2; end
			4413: begin bcd3<=4;bcd2<=4;bcd1<=1;bcd0<=3; end
			4414: begin bcd3<=4;bcd2<=4;bcd1<=1;bcd0<=4; end
			4415: begin bcd3<=4;bcd2<=4;bcd1<=1;bcd0<=5; end
			4416: begin bcd3<=4;bcd2<=4;bcd1<=1;bcd0<=6; end
			4417: begin bcd3<=4;bcd2<=4;bcd1<=1;bcd0<=7; end
			4418: begin bcd3<=4;bcd2<=4;bcd1<=1;bcd0<=8; end
			4419: begin bcd3<=4;bcd2<=4;bcd1<=1;bcd0<=9; end
			4420: begin bcd3<=4;bcd2<=4;bcd1<=2;bcd0<=0; end
			4421: begin bcd3<=4;bcd2<=4;bcd1<=2;bcd0<=1; end
			4422: begin bcd3<=4;bcd2<=4;bcd1<=2;bcd0<=2; end
			4423: begin bcd3<=4;bcd2<=4;bcd1<=2;bcd0<=3; end
			4424: begin bcd3<=4;bcd2<=4;bcd1<=2;bcd0<=4; end
			4425: begin bcd3<=4;bcd2<=4;bcd1<=2;bcd0<=5; end
			4426: begin bcd3<=4;bcd2<=4;bcd1<=2;bcd0<=6; end
			4427: begin bcd3<=4;bcd2<=4;bcd1<=2;bcd0<=7; end
			4428: begin bcd3<=4;bcd2<=4;bcd1<=2;bcd0<=8; end
			4429: begin bcd3<=4;bcd2<=4;bcd1<=2;bcd0<=9; end
			4430: begin bcd3<=4;bcd2<=4;bcd1<=3;bcd0<=0; end
			4431: begin bcd3<=4;bcd2<=4;bcd1<=3;bcd0<=1; end
			4432: begin bcd3<=4;bcd2<=4;bcd1<=3;bcd0<=2; end
			4433: begin bcd3<=4;bcd2<=4;bcd1<=3;bcd0<=3; end
			4434: begin bcd3<=4;bcd2<=4;bcd1<=3;bcd0<=4; end
			4435: begin bcd3<=4;bcd2<=4;bcd1<=3;bcd0<=5; end
			4436: begin bcd3<=4;bcd2<=4;bcd1<=3;bcd0<=6; end
			4437: begin bcd3<=4;bcd2<=4;bcd1<=3;bcd0<=7; end
			4438: begin bcd3<=4;bcd2<=4;bcd1<=3;bcd0<=8; end
			4439: begin bcd3<=4;bcd2<=4;bcd1<=3;bcd0<=9; end
			4440: begin bcd3<=4;bcd2<=4;bcd1<=4;bcd0<=0; end
			4441: begin bcd3<=4;bcd2<=4;bcd1<=4;bcd0<=1; end
			4442: begin bcd3<=4;bcd2<=4;bcd1<=4;bcd0<=2; end
			4443: begin bcd3<=4;bcd2<=4;bcd1<=4;bcd0<=3; end
			4444: begin bcd3<=4;bcd2<=4;bcd1<=4;bcd0<=4; end
			4445: begin bcd3<=4;bcd2<=4;bcd1<=4;bcd0<=5; end
			4446: begin bcd3<=4;bcd2<=4;bcd1<=4;bcd0<=6; end
			4447: begin bcd3<=4;bcd2<=4;bcd1<=4;bcd0<=7; end
			4448: begin bcd3<=4;bcd2<=4;bcd1<=4;bcd0<=8; end
			4449: begin bcd3<=4;bcd2<=4;bcd1<=4;bcd0<=9; end
			4450: begin bcd3<=4;bcd2<=4;bcd1<=5;bcd0<=0; end
			4451: begin bcd3<=4;bcd2<=4;bcd1<=5;bcd0<=1; end
			4452: begin bcd3<=4;bcd2<=4;bcd1<=5;bcd0<=2; end
			4453: begin bcd3<=4;bcd2<=4;bcd1<=5;bcd0<=3; end
			4454: begin bcd3<=4;bcd2<=4;bcd1<=5;bcd0<=4; end
			4455: begin bcd3<=4;bcd2<=4;bcd1<=5;bcd0<=5; end
			4456: begin bcd3<=4;bcd2<=4;bcd1<=5;bcd0<=6; end
			4457: begin bcd3<=4;bcd2<=4;bcd1<=5;bcd0<=7; end
			4458: begin bcd3<=4;bcd2<=4;bcd1<=5;bcd0<=8; end
			4459: begin bcd3<=4;bcd2<=4;bcd1<=5;bcd0<=9; end
			4460: begin bcd3<=4;bcd2<=4;bcd1<=6;bcd0<=0; end
			4461: begin bcd3<=4;bcd2<=4;bcd1<=6;bcd0<=1; end
			4462: begin bcd3<=4;bcd2<=4;bcd1<=6;bcd0<=2; end
			4463: begin bcd3<=4;bcd2<=4;bcd1<=6;bcd0<=3; end
			4464: begin bcd3<=4;bcd2<=4;bcd1<=6;bcd0<=4; end
			4465: begin bcd3<=4;bcd2<=4;bcd1<=6;bcd0<=5; end
			4466: begin bcd3<=4;bcd2<=4;bcd1<=6;bcd0<=6; end
			4467: begin bcd3<=4;bcd2<=4;bcd1<=6;bcd0<=7; end
			4468: begin bcd3<=4;bcd2<=4;bcd1<=6;bcd0<=8; end
			4469: begin bcd3<=4;bcd2<=4;bcd1<=6;bcd0<=9; end
			4470: begin bcd3<=4;bcd2<=4;bcd1<=7;bcd0<=0; end
			4471: begin bcd3<=4;bcd2<=4;bcd1<=7;bcd0<=1; end
			4472: begin bcd3<=4;bcd2<=4;bcd1<=7;bcd0<=2; end
			4473: begin bcd3<=4;bcd2<=4;bcd1<=7;bcd0<=3; end
			4474: begin bcd3<=4;bcd2<=4;bcd1<=7;bcd0<=4; end
			4475: begin bcd3<=4;bcd2<=4;bcd1<=7;bcd0<=5; end
			4476: begin bcd3<=4;bcd2<=4;bcd1<=7;bcd0<=6; end
			4477: begin bcd3<=4;bcd2<=4;bcd1<=7;bcd0<=7; end
			4478: begin bcd3<=4;bcd2<=4;bcd1<=7;bcd0<=8; end
			4479: begin bcd3<=4;bcd2<=4;bcd1<=7;bcd0<=9; end
			4480: begin bcd3<=4;bcd2<=4;bcd1<=8;bcd0<=0; end
			4481: begin bcd3<=4;bcd2<=4;bcd1<=8;bcd0<=1; end
			4482: begin bcd3<=4;bcd2<=4;bcd1<=8;bcd0<=2; end
			4483: begin bcd3<=4;bcd2<=4;bcd1<=8;bcd0<=3; end
			4484: begin bcd3<=4;bcd2<=4;bcd1<=8;bcd0<=4; end
			4485: begin bcd3<=4;bcd2<=4;bcd1<=8;bcd0<=5; end
			4486: begin bcd3<=4;bcd2<=4;bcd1<=8;bcd0<=6; end
			4487: begin bcd3<=4;bcd2<=4;bcd1<=8;bcd0<=7; end
			4488: begin bcd3<=4;bcd2<=4;bcd1<=8;bcd0<=8; end
			4489: begin bcd3<=4;bcd2<=4;bcd1<=8;bcd0<=9; end
			4490: begin bcd3<=4;bcd2<=4;bcd1<=9;bcd0<=0; end
			4491: begin bcd3<=4;bcd2<=4;bcd1<=9;bcd0<=1; end
			4492: begin bcd3<=4;bcd2<=4;bcd1<=9;bcd0<=2; end
			4493: begin bcd3<=4;bcd2<=4;bcd1<=9;bcd0<=3; end
			4494: begin bcd3<=4;bcd2<=4;bcd1<=9;bcd0<=4; end
			4495: begin bcd3<=4;bcd2<=4;bcd1<=9;bcd0<=5; end
			4496: begin bcd3<=4;bcd2<=4;bcd1<=9;bcd0<=6; end
			4497: begin bcd3<=4;bcd2<=4;bcd1<=9;bcd0<=7; end
			4498: begin bcd3<=4;bcd2<=4;bcd1<=9;bcd0<=8; end
			4499: begin bcd3<=4;bcd2<=4;bcd1<=9;bcd0<=9; end
			4500: begin bcd3<=4;bcd2<=5;bcd1<=0;bcd0<=0; end
			4501: begin bcd3<=4;bcd2<=5;bcd1<=0;bcd0<=1; end
			4502: begin bcd3<=4;bcd2<=5;bcd1<=0;bcd0<=2; end
			4503: begin bcd3<=4;bcd2<=5;bcd1<=0;bcd0<=3; end
			4504: begin bcd3<=4;bcd2<=5;bcd1<=0;bcd0<=4; end
			4505: begin bcd3<=4;bcd2<=5;bcd1<=0;bcd0<=5; end
			4506: begin bcd3<=4;bcd2<=5;bcd1<=0;bcd0<=6; end
			4507: begin bcd3<=4;bcd2<=5;bcd1<=0;bcd0<=7; end
			4508: begin bcd3<=4;bcd2<=5;bcd1<=0;bcd0<=8; end
			4509: begin bcd3<=4;bcd2<=5;bcd1<=0;bcd0<=9; end
			4510: begin bcd3<=4;bcd2<=5;bcd1<=1;bcd0<=0; end
			4511: begin bcd3<=4;bcd2<=5;bcd1<=1;bcd0<=1; end
			4512: begin bcd3<=4;bcd2<=5;bcd1<=1;bcd0<=2; end
			4513: begin bcd3<=4;bcd2<=5;bcd1<=1;bcd0<=3; end
			4514: begin bcd3<=4;bcd2<=5;bcd1<=1;bcd0<=4; end
			4515: begin bcd3<=4;bcd2<=5;bcd1<=1;bcd0<=5; end
			4516: begin bcd3<=4;bcd2<=5;bcd1<=1;bcd0<=6; end
			4517: begin bcd3<=4;bcd2<=5;bcd1<=1;bcd0<=7; end
			4518: begin bcd3<=4;bcd2<=5;bcd1<=1;bcd0<=8; end
			4519: begin bcd3<=4;bcd2<=5;bcd1<=1;bcd0<=9; end
			4520: begin bcd3<=4;bcd2<=5;bcd1<=2;bcd0<=0; end
			4521: begin bcd3<=4;bcd2<=5;bcd1<=2;bcd0<=1; end
			4522: begin bcd3<=4;bcd2<=5;bcd1<=2;bcd0<=2; end
			4523: begin bcd3<=4;bcd2<=5;bcd1<=2;bcd0<=3; end
			4524: begin bcd3<=4;bcd2<=5;bcd1<=2;bcd0<=4; end
			4525: begin bcd3<=4;bcd2<=5;bcd1<=2;bcd0<=5; end
			4526: begin bcd3<=4;bcd2<=5;bcd1<=2;bcd0<=6; end
			4527: begin bcd3<=4;bcd2<=5;bcd1<=2;bcd0<=7; end
			4528: begin bcd3<=4;bcd2<=5;bcd1<=2;bcd0<=8; end
			4529: begin bcd3<=4;bcd2<=5;bcd1<=2;bcd0<=9; end
			4530: begin bcd3<=4;bcd2<=5;bcd1<=3;bcd0<=0; end
			4531: begin bcd3<=4;bcd2<=5;bcd1<=3;bcd0<=1; end
			4532: begin bcd3<=4;bcd2<=5;bcd1<=3;bcd0<=2; end
			4533: begin bcd3<=4;bcd2<=5;bcd1<=3;bcd0<=3; end
			4534: begin bcd3<=4;bcd2<=5;bcd1<=3;bcd0<=4; end
			4535: begin bcd3<=4;bcd2<=5;bcd1<=3;bcd0<=5; end
			4536: begin bcd3<=4;bcd2<=5;bcd1<=3;bcd0<=6; end
			4537: begin bcd3<=4;bcd2<=5;bcd1<=3;bcd0<=7; end
			4538: begin bcd3<=4;bcd2<=5;bcd1<=3;bcd0<=8; end
			4539: begin bcd3<=4;bcd2<=5;bcd1<=3;bcd0<=9; end
			4540: begin bcd3<=4;bcd2<=5;bcd1<=4;bcd0<=0; end
			4541: begin bcd3<=4;bcd2<=5;bcd1<=4;bcd0<=1; end
			4542: begin bcd3<=4;bcd2<=5;bcd1<=4;bcd0<=2; end
			4543: begin bcd3<=4;bcd2<=5;bcd1<=4;bcd0<=3; end
			4544: begin bcd3<=4;bcd2<=5;bcd1<=4;bcd0<=4; end
			4545: begin bcd3<=4;bcd2<=5;bcd1<=4;bcd0<=5; end
			4546: begin bcd3<=4;bcd2<=5;bcd1<=4;bcd0<=6; end
			4547: begin bcd3<=4;bcd2<=5;bcd1<=4;bcd0<=7; end
			4548: begin bcd3<=4;bcd2<=5;bcd1<=4;bcd0<=8; end
			4549: begin bcd3<=4;bcd2<=5;bcd1<=4;bcd0<=9; end
			4550: begin bcd3<=4;bcd2<=5;bcd1<=5;bcd0<=0; end
			4551: begin bcd3<=4;bcd2<=5;bcd1<=5;bcd0<=1; end
			4552: begin bcd3<=4;bcd2<=5;bcd1<=5;bcd0<=2; end
			4553: begin bcd3<=4;bcd2<=5;bcd1<=5;bcd0<=3; end
			4554: begin bcd3<=4;bcd2<=5;bcd1<=5;bcd0<=4; end
			4555: begin bcd3<=4;bcd2<=5;bcd1<=5;bcd0<=5; end
			4556: begin bcd3<=4;bcd2<=5;bcd1<=5;bcd0<=6; end
			4557: begin bcd3<=4;bcd2<=5;bcd1<=5;bcd0<=7; end
			4558: begin bcd3<=4;bcd2<=5;bcd1<=5;bcd0<=8; end
			4559: begin bcd3<=4;bcd2<=5;bcd1<=5;bcd0<=9; end
			4560: begin bcd3<=4;bcd2<=5;bcd1<=6;bcd0<=0; end
			4561: begin bcd3<=4;bcd2<=5;bcd1<=6;bcd0<=1; end
			4562: begin bcd3<=4;bcd2<=5;bcd1<=6;bcd0<=2; end
			4563: begin bcd3<=4;bcd2<=5;bcd1<=6;bcd0<=3; end
			4564: begin bcd3<=4;bcd2<=5;bcd1<=6;bcd0<=4; end
			4565: begin bcd3<=4;bcd2<=5;bcd1<=6;bcd0<=5; end
			4566: begin bcd3<=4;bcd2<=5;bcd1<=6;bcd0<=6; end
			4567: begin bcd3<=4;bcd2<=5;bcd1<=6;bcd0<=7; end
			4568: begin bcd3<=4;bcd2<=5;bcd1<=6;bcd0<=8; end
			4569: begin bcd3<=4;bcd2<=5;bcd1<=6;bcd0<=9; end
			4570: begin bcd3<=4;bcd2<=5;bcd1<=7;bcd0<=0; end
			4571: begin bcd3<=4;bcd2<=5;bcd1<=7;bcd0<=1; end
			4572: begin bcd3<=4;bcd2<=5;bcd1<=7;bcd0<=2; end
			4573: begin bcd3<=4;bcd2<=5;bcd1<=7;bcd0<=3; end
			4574: begin bcd3<=4;bcd2<=5;bcd1<=7;bcd0<=4; end
			4575: begin bcd3<=4;bcd2<=5;bcd1<=7;bcd0<=5; end
			4576: begin bcd3<=4;bcd2<=5;bcd1<=7;bcd0<=6; end
			4577: begin bcd3<=4;bcd2<=5;bcd1<=7;bcd0<=7; end
			4578: begin bcd3<=4;bcd2<=5;bcd1<=7;bcd0<=8; end
			4579: begin bcd3<=4;bcd2<=5;bcd1<=7;bcd0<=9; end
			4580: begin bcd3<=4;bcd2<=5;bcd1<=8;bcd0<=0; end
			4581: begin bcd3<=4;bcd2<=5;bcd1<=8;bcd0<=1; end
			4582: begin bcd3<=4;bcd2<=5;bcd1<=8;bcd0<=2; end
			4583: begin bcd3<=4;bcd2<=5;bcd1<=8;bcd0<=3; end
			4584: begin bcd3<=4;bcd2<=5;bcd1<=8;bcd0<=4; end
			4585: begin bcd3<=4;bcd2<=5;bcd1<=8;bcd0<=5; end
			4586: begin bcd3<=4;bcd2<=5;bcd1<=8;bcd0<=6; end
			4587: begin bcd3<=4;bcd2<=5;bcd1<=8;bcd0<=7; end
			4588: begin bcd3<=4;bcd2<=5;bcd1<=8;bcd0<=8; end
			4589: begin bcd3<=4;bcd2<=5;bcd1<=8;bcd0<=9; end
			4590: begin bcd3<=4;bcd2<=5;bcd1<=9;bcd0<=0; end
			4591: begin bcd3<=4;bcd2<=5;bcd1<=9;bcd0<=1; end
			4592: begin bcd3<=4;bcd2<=5;bcd1<=9;bcd0<=2; end
			4593: begin bcd3<=4;bcd2<=5;bcd1<=9;bcd0<=3; end
			4594: begin bcd3<=4;bcd2<=5;bcd1<=9;bcd0<=4; end
			4595: begin bcd3<=4;bcd2<=5;bcd1<=9;bcd0<=5; end
			4596: begin bcd3<=4;bcd2<=5;bcd1<=9;bcd0<=6; end
			4597: begin bcd3<=4;bcd2<=5;bcd1<=9;bcd0<=7; end
			4598: begin bcd3<=4;bcd2<=5;bcd1<=9;bcd0<=8; end
			4599: begin bcd3<=4;bcd2<=5;bcd1<=9;bcd0<=9; end
			4600: begin bcd3<=4;bcd2<=6;bcd1<=0;bcd0<=0; end
			4601: begin bcd3<=4;bcd2<=6;bcd1<=0;bcd0<=1; end
			4602: begin bcd3<=4;bcd2<=6;bcd1<=0;bcd0<=2; end
			4603: begin bcd3<=4;bcd2<=6;bcd1<=0;bcd0<=3; end
			4604: begin bcd3<=4;bcd2<=6;bcd1<=0;bcd0<=4; end
			4605: begin bcd3<=4;bcd2<=6;bcd1<=0;bcd0<=5; end
			4606: begin bcd3<=4;bcd2<=6;bcd1<=0;bcd0<=6; end
			4607: begin bcd3<=4;bcd2<=6;bcd1<=0;bcd0<=7; end
			4608: begin bcd3<=4;bcd2<=6;bcd1<=0;bcd0<=8; end
			4609: begin bcd3<=4;bcd2<=6;bcd1<=0;bcd0<=9; end
			4610: begin bcd3<=4;bcd2<=6;bcd1<=1;bcd0<=0; end
			4611: begin bcd3<=4;bcd2<=6;bcd1<=1;bcd0<=1; end
			4612: begin bcd3<=4;bcd2<=6;bcd1<=1;bcd0<=2; end
			4613: begin bcd3<=4;bcd2<=6;bcd1<=1;bcd0<=3; end
			4614: begin bcd3<=4;bcd2<=6;bcd1<=1;bcd0<=4; end
			4615: begin bcd3<=4;bcd2<=6;bcd1<=1;bcd0<=5; end
			4616: begin bcd3<=4;bcd2<=6;bcd1<=1;bcd0<=6; end
			4617: begin bcd3<=4;bcd2<=6;bcd1<=1;bcd0<=7; end
			4618: begin bcd3<=4;bcd2<=6;bcd1<=1;bcd0<=8; end
			4619: begin bcd3<=4;bcd2<=6;bcd1<=1;bcd0<=9; end
			4620: begin bcd3<=4;bcd2<=6;bcd1<=2;bcd0<=0; end
			4621: begin bcd3<=4;bcd2<=6;bcd1<=2;bcd0<=1; end
			4622: begin bcd3<=4;bcd2<=6;bcd1<=2;bcd0<=2; end
			4623: begin bcd3<=4;bcd2<=6;bcd1<=2;bcd0<=3; end
			4624: begin bcd3<=4;bcd2<=6;bcd1<=2;bcd0<=4; end
			4625: begin bcd3<=4;bcd2<=6;bcd1<=2;bcd0<=5; end
			4626: begin bcd3<=4;bcd2<=6;bcd1<=2;bcd0<=6; end
			4627: begin bcd3<=4;bcd2<=6;bcd1<=2;bcd0<=7; end
			4628: begin bcd3<=4;bcd2<=6;bcd1<=2;bcd0<=8; end
			4629: begin bcd3<=4;bcd2<=6;bcd1<=2;bcd0<=9; end
			4630: begin bcd3<=4;bcd2<=6;bcd1<=3;bcd0<=0; end
			4631: begin bcd3<=4;bcd2<=6;bcd1<=3;bcd0<=1; end
			4632: begin bcd3<=4;bcd2<=6;bcd1<=3;bcd0<=2; end
			4633: begin bcd3<=4;bcd2<=6;bcd1<=3;bcd0<=3; end
			4634: begin bcd3<=4;bcd2<=6;bcd1<=3;bcd0<=4; end
			4635: begin bcd3<=4;bcd2<=6;bcd1<=3;bcd0<=5; end
			4636: begin bcd3<=4;bcd2<=6;bcd1<=3;bcd0<=6; end
			4637: begin bcd3<=4;bcd2<=6;bcd1<=3;bcd0<=7; end
			4638: begin bcd3<=4;bcd2<=6;bcd1<=3;bcd0<=8; end
			4639: begin bcd3<=4;bcd2<=6;bcd1<=3;bcd0<=9; end
			4640: begin bcd3<=4;bcd2<=6;bcd1<=4;bcd0<=0; end
			4641: begin bcd3<=4;bcd2<=6;bcd1<=4;bcd0<=1; end
			4642: begin bcd3<=4;bcd2<=6;bcd1<=4;bcd0<=2; end
			4643: begin bcd3<=4;bcd2<=6;bcd1<=4;bcd0<=3; end
			4644: begin bcd3<=4;bcd2<=6;bcd1<=4;bcd0<=4; end
			4645: begin bcd3<=4;bcd2<=6;bcd1<=4;bcd0<=5; end
			4646: begin bcd3<=4;bcd2<=6;bcd1<=4;bcd0<=6; end
			4647: begin bcd3<=4;bcd2<=6;bcd1<=4;bcd0<=7; end
			4648: begin bcd3<=4;bcd2<=6;bcd1<=4;bcd0<=8; end
			4649: begin bcd3<=4;bcd2<=6;bcd1<=4;bcd0<=9; end
			4650: begin bcd3<=4;bcd2<=6;bcd1<=5;bcd0<=0; end
			4651: begin bcd3<=4;bcd2<=6;bcd1<=5;bcd0<=1; end
			4652: begin bcd3<=4;bcd2<=6;bcd1<=5;bcd0<=2; end
			4653: begin bcd3<=4;bcd2<=6;bcd1<=5;bcd0<=3; end
			4654: begin bcd3<=4;bcd2<=6;bcd1<=5;bcd0<=4; end
			4655: begin bcd3<=4;bcd2<=6;bcd1<=5;bcd0<=5; end
			4656: begin bcd3<=4;bcd2<=6;bcd1<=5;bcd0<=6; end
			4657: begin bcd3<=4;bcd2<=6;bcd1<=5;bcd0<=7; end
			4658: begin bcd3<=4;bcd2<=6;bcd1<=5;bcd0<=8; end
			4659: begin bcd3<=4;bcd2<=6;bcd1<=5;bcd0<=9; end
			4660: begin bcd3<=4;bcd2<=6;bcd1<=6;bcd0<=0; end
			4661: begin bcd3<=4;bcd2<=6;bcd1<=6;bcd0<=1; end
			4662: begin bcd3<=4;bcd2<=6;bcd1<=6;bcd0<=2; end
			4663: begin bcd3<=4;bcd2<=6;bcd1<=6;bcd0<=3; end
			4664: begin bcd3<=4;bcd2<=6;bcd1<=6;bcd0<=4; end
			4665: begin bcd3<=4;bcd2<=6;bcd1<=6;bcd0<=5; end
			4666: begin bcd3<=4;bcd2<=6;bcd1<=6;bcd0<=6; end
			4667: begin bcd3<=4;bcd2<=6;bcd1<=6;bcd0<=7; end
			4668: begin bcd3<=4;bcd2<=6;bcd1<=6;bcd0<=8; end
			4669: begin bcd3<=4;bcd2<=6;bcd1<=6;bcd0<=9; end
			4670: begin bcd3<=4;bcd2<=6;bcd1<=7;bcd0<=0; end
			4671: begin bcd3<=4;bcd2<=6;bcd1<=7;bcd0<=1; end
			4672: begin bcd3<=4;bcd2<=6;bcd1<=7;bcd0<=2; end
			4673: begin bcd3<=4;bcd2<=6;bcd1<=7;bcd0<=3; end
			4674: begin bcd3<=4;bcd2<=6;bcd1<=7;bcd0<=4; end
			4675: begin bcd3<=4;bcd2<=6;bcd1<=7;bcd0<=5; end
			4676: begin bcd3<=4;bcd2<=6;bcd1<=7;bcd0<=6; end
			4677: begin bcd3<=4;bcd2<=6;bcd1<=7;bcd0<=7; end
			4678: begin bcd3<=4;bcd2<=6;bcd1<=7;bcd0<=8; end
			4679: begin bcd3<=4;bcd2<=6;bcd1<=7;bcd0<=9; end
			4680: begin bcd3<=4;bcd2<=6;bcd1<=8;bcd0<=0; end
			4681: begin bcd3<=4;bcd2<=6;bcd1<=8;bcd0<=1; end
			4682: begin bcd3<=4;bcd2<=6;bcd1<=8;bcd0<=2; end
			4683: begin bcd3<=4;bcd2<=6;bcd1<=8;bcd0<=3; end
			4684: begin bcd3<=4;bcd2<=6;bcd1<=8;bcd0<=4; end
			4685: begin bcd3<=4;bcd2<=6;bcd1<=8;bcd0<=5; end
			4686: begin bcd3<=4;bcd2<=6;bcd1<=8;bcd0<=6; end
			4687: begin bcd3<=4;bcd2<=6;bcd1<=8;bcd0<=7; end
			4688: begin bcd3<=4;bcd2<=6;bcd1<=8;bcd0<=8; end
			4689: begin bcd3<=4;bcd2<=6;bcd1<=8;bcd0<=9; end
			4690: begin bcd3<=4;bcd2<=6;bcd1<=9;bcd0<=0; end
			4691: begin bcd3<=4;bcd2<=6;bcd1<=9;bcd0<=1; end
			4692: begin bcd3<=4;bcd2<=6;bcd1<=9;bcd0<=2; end
			4693: begin bcd3<=4;bcd2<=6;bcd1<=9;bcd0<=3; end
			4694: begin bcd3<=4;bcd2<=6;bcd1<=9;bcd0<=4; end
			4695: begin bcd3<=4;bcd2<=6;bcd1<=9;bcd0<=5; end
			4696: begin bcd3<=4;bcd2<=6;bcd1<=9;bcd0<=6; end
			4697: begin bcd3<=4;bcd2<=6;bcd1<=9;bcd0<=7; end
			4698: begin bcd3<=4;bcd2<=6;bcd1<=9;bcd0<=8; end
			4699: begin bcd3<=4;bcd2<=6;bcd1<=9;bcd0<=9; end
			4700: begin bcd3<=4;bcd2<=7;bcd1<=0;bcd0<=0; end
			4701: begin bcd3<=4;bcd2<=7;bcd1<=0;bcd0<=1; end
			4702: begin bcd3<=4;bcd2<=7;bcd1<=0;bcd0<=2; end
			4703: begin bcd3<=4;bcd2<=7;bcd1<=0;bcd0<=3; end
			4704: begin bcd3<=4;bcd2<=7;bcd1<=0;bcd0<=4; end
			4705: begin bcd3<=4;bcd2<=7;bcd1<=0;bcd0<=5; end
			4706: begin bcd3<=4;bcd2<=7;bcd1<=0;bcd0<=6; end
			4707: begin bcd3<=4;bcd2<=7;bcd1<=0;bcd0<=7; end
			4708: begin bcd3<=4;bcd2<=7;bcd1<=0;bcd0<=8; end
			4709: begin bcd3<=4;bcd2<=7;bcd1<=0;bcd0<=9; end
			4710: begin bcd3<=4;bcd2<=7;bcd1<=1;bcd0<=0; end
			4711: begin bcd3<=4;bcd2<=7;bcd1<=1;bcd0<=1; end
			4712: begin bcd3<=4;bcd2<=7;bcd1<=1;bcd0<=2; end
			4713: begin bcd3<=4;bcd2<=7;bcd1<=1;bcd0<=3; end
			4714: begin bcd3<=4;bcd2<=7;bcd1<=1;bcd0<=4; end
			4715: begin bcd3<=4;bcd2<=7;bcd1<=1;bcd0<=5; end
			4716: begin bcd3<=4;bcd2<=7;bcd1<=1;bcd0<=6; end
			4717: begin bcd3<=4;bcd2<=7;bcd1<=1;bcd0<=7; end
			4718: begin bcd3<=4;bcd2<=7;bcd1<=1;bcd0<=8; end
			4719: begin bcd3<=4;bcd2<=7;bcd1<=1;bcd0<=9; end
			4720: begin bcd3<=4;bcd2<=7;bcd1<=2;bcd0<=0; end
			4721: begin bcd3<=4;bcd2<=7;bcd1<=2;bcd0<=1; end
			4722: begin bcd3<=4;bcd2<=7;bcd1<=2;bcd0<=2; end
			4723: begin bcd3<=4;bcd2<=7;bcd1<=2;bcd0<=3; end
			4724: begin bcd3<=4;bcd2<=7;bcd1<=2;bcd0<=4; end
			4725: begin bcd3<=4;bcd2<=7;bcd1<=2;bcd0<=5; end
			4726: begin bcd3<=4;bcd2<=7;bcd1<=2;bcd0<=6; end
			4727: begin bcd3<=4;bcd2<=7;bcd1<=2;bcd0<=7; end
			4728: begin bcd3<=4;bcd2<=7;bcd1<=2;bcd0<=8; end
			4729: begin bcd3<=4;bcd2<=7;bcd1<=2;bcd0<=9; end
			4730: begin bcd3<=4;bcd2<=7;bcd1<=3;bcd0<=0; end
			4731: begin bcd3<=4;bcd2<=7;bcd1<=3;bcd0<=1; end
			4732: begin bcd3<=4;bcd2<=7;bcd1<=3;bcd0<=2; end
			4733: begin bcd3<=4;bcd2<=7;bcd1<=3;bcd0<=3; end
			4734: begin bcd3<=4;bcd2<=7;bcd1<=3;bcd0<=4; end
			4735: begin bcd3<=4;bcd2<=7;bcd1<=3;bcd0<=5; end
			4736: begin bcd3<=4;bcd2<=7;bcd1<=3;bcd0<=6; end
			4737: begin bcd3<=4;bcd2<=7;bcd1<=3;bcd0<=7; end
			4738: begin bcd3<=4;bcd2<=7;bcd1<=3;bcd0<=8; end
			4739: begin bcd3<=4;bcd2<=7;bcd1<=3;bcd0<=9; end
			4740: begin bcd3<=4;bcd2<=7;bcd1<=4;bcd0<=0; end
			4741: begin bcd3<=4;bcd2<=7;bcd1<=4;bcd0<=1; end
			4742: begin bcd3<=4;bcd2<=7;bcd1<=4;bcd0<=2; end
			4743: begin bcd3<=4;bcd2<=7;bcd1<=4;bcd0<=3; end
			4744: begin bcd3<=4;bcd2<=7;bcd1<=4;bcd0<=4; end
			4745: begin bcd3<=4;bcd2<=7;bcd1<=4;bcd0<=5; end
			4746: begin bcd3<=4;bcd2<=7;bcd1<=4;bcd0<=6; end
			4747: begin bcd3<=4;bcd2<=7;bcd1<=4;bcd0<=7; end
			4748: begin bcd3<=4;bcd2<=7;bcd1<=4;bcd0<=8; end
			4749: begin bcd3<=4;bcd2<=7;bcd1<=4;bcd0<=9; end
			4750: begin bcd3<=4;bcd2<=7;bcd1<=5;bcd0<=0; end
			4751: begin bcd3<=4;bcd2<=7;bcd1<=5;bcd0<=1; end
			4752: begin bcd3<=4;bcd2<=7;bcd1<=5;bcd0<=2; end
			4753: begin bcd3<=4;bcd2<=7;bcd1<=5;bcd0<=3; end
			4754: begin bcd3<=4;bcd2<=7;bcd1<=5;bcd0<=4; end
			4755: begin bcd3<=4;bcd2<=7;bcd1<=5;bcd0<=5; end
			4756: begin bcd3<=4;bcd2<=7;bcd1<=5;bcd0<=6; end
			4757: begin bcd3<=4;bcd2<=7;bcd1<=5;bcd0<=7; end
			4758: begin bcd3<=4;bcd2<=7;bcd1<=5;bcd0<=8; end
			4759: begin bcd3<=4;bcd2<=7;bcd1<=5;bcd0<=9; end
			4760: begin bcd3<=4;bcd2<=7;bcd1<=6;bcd0<=0; end
			4761: begin bcd3<=4;bcd2<=7;bcd1<=6;bcd0<=1; end
			4762: begin bcd3<=4;bcd2<=7;bcd1<=6;bcd0<=2; end
			4763: begin bcd3<=4;bcd2<=7;bcd1<=6;bcd0<=3; end
			4764: begin bcd3<=4;bcd2<=7;bcd1<=6;bcd0<=4; end
			4765: begin bcd3<=4;bcd2<=7;bcd1<=6;bcd0<=5; end
			4766: begin bcd3<=4;bcd2<=7;bcd1<=6;bcd0<=6; end
			4767: begin bcd3<=4;bcd2<=7;bcd1<=6;bcd0<=7; end
			4768: begin bcd3<=4;bcd2<=7;bcd1<=6;bcd0<=8; end
			4769: begin bcd3<=4;bcd2<=7;bcd1<=6;bcd0<=9; end
			4770: begin bcd3<=4;bcd2<=7;bcd1<=7;bcd0<=0; end
			4771: begin bcd3<=4;bcd2<=7;bcd1<=7;bcd0<=1; end
			4772: begin bcd3<=4;bcd2<=7;bcd1<=7;bcd0<=2; end
			4773: begin bcd3<=4;bcd2<=7;bcd1<=7;bcd0<=3; end
			4774: begin bcd3<=4;bcd2<=7;bcd1<=7;bcd0<=4; end
			4775: begin bcd3<=4;bcd2<=7;bcd1<=7;bcd0<=5; end
			4776: begin bcd3<=4;bcd2<=7;bcd1<=7;bcd0<=6; end
			4777: begin bcd3<=4;bcd2<=7;bcd1<=7;bcd0<=7; end
			4778: begin bcd3<=4;bcd2<=7;bcd1<=7;bcd0<=8; end
			4779: begin bcd3<=4;bcd2<=7;bcd1<=7;bcd0<=9; end
			4780: begin bcd3<=4;bcd2<=7;bcd1<=8;bcd0<=0; end
			4781: begin bcd3<=4;bcd2<=7;bcd1<=8;bcd0<=1; end
			4782: begin bcd3<=4;bcd2<=7;bcd1<=8;bcd0<=2; end
			4783: begin bcd3<=4;bcd2<=7;bcd1<=8;bcd0<=3; end
			4784: begin bcd3<=4;bcd2<=7;bcd1<=8;bcd0<=4; end
			4785: begin bcd3<=4;bcd2<=7;bcd1<=8;bcd0<=5; end
			4786: begin bcd3<=4;bcd2<=7;bcd1<=8;bcd0<=6; end
			4787: begin bcd3<=4;bcd2<=7;bcd1<=8;bcd0<=7; end
			4788: begin bcd3<=4;bcd2<=7;bcd1<=8;bcd0<=8; end
			4789: begin bcd3<=4;bcd2<=7;bcd1<=8;bcd0<=9; end
			4790: begin bcd3<=4;bcd2<=7;bcd1<=9;bcd0<=0; end
			4791: begin bcd3<=4;bcd2<=7;bcd1<=9;bcd0<=1; end
			4792: begin bcd3<=4;bcd2<=7;bcd1<=9;bcd0<=2; end
			4793: begin bcd3<=4;bcd2<=7;bcd1<=9;bcd0<=3; end
			4794: begin bcd3<=4;bcd2<=7;bcd1<=9;bcd0<=4; end
			4795: begin bcd3<=4;bcd2<=7;bcd1<=9;bcd0<=5; end
			4796: begin bcd3<=4;bcd2<=7;bcd1<=9;bcd0<=6; end
			4797: begin bcd3<=4;bcd2<=7;bcd1<=9;bcd0<=7; end
			4798: begin bcd3<=4;bcd2<=7;bcd1<=9;bcd0<=8; end
			4799: begin bcd3<=4;bcd2<=7;bcd1<=9;bcd0<=9; end
			4800: begin bcd3<=4;bcd2<=8;bcd1<=0;bcd0<=0; end
			4801: begin bcd3<=4;bcd2<=8;bcd1<=0;bcd0<=1; end
			4802: begin bcd3<=4;bcd2<=8;bcd1<=0;bcd0<=2; end
			4803: begin bcd3<=4;bcd2<=8;bcd1<=0;bcd0<=3; end
			4804: begin bcd3<=4;bcd2<=8;bcd1<=0;bcd0<=4; end
			4805: begin bcd3<=4;bcd2<=8;bcd1<=0;bcd0<=5; end
			4806: begin bcd3<=4;bcd2<=8;bcd1<=0;bcd0<=6; end
			4807: begin bcd3<=4;bcd2<=8;bcd1<=0;bcd0<=7; end
			4808: begin bcd3<=4;bcd2<=8;bcd1<=0;bcd0<=8; end
			4809: begin bcd3<=4;bcd2<=8;bcd1<=0;bcd0<=9; end
			4810: begin bcd3<=4;bcd2<=8;bcd1<=1;bcd0<=0; end
			4811: begin bcd3<=4;bcd2<=8;bcd1<=1;bcd0<=1; end
			4812: begin bcd3<=4;bcd2<=8;bcd1<=1;bcd0<=2; end
			4813: begin bcd3<=4;bcd2<=8;bcd1<=1;bcd0<=3; end
			4814: begin bcd3<=4;bcd2<=8;bcd1<=1;bcd0<=4; end
			4815: begin bcd3<=4;bcd2<=8;bcd1<=1;bcd0<=5; end
			4816: begin bcd3<=4;bcd2<=8;bcd1<=1;bcd0<=6; end
			4817: begin bcd3<=4;bcd2<=8;bcd1<=1;bcd0<=7; end
			4818: begin bcd3<=4;bcd2<=8;bcd1<=1;bcd0<=8; end
			4819: begin bcd3<=4;bcd2<=8;bcd1<=1;bcd0<=9; end
			4820: begin bcd3<=4;bcd2<=8;bcd1<=2;bcd0<=0; end
			4821: begin bcd3<=4;bcd2<=8;bcd1<=2;bcd0<=1; end
			4822: begin bcd3<=4;bcd2<=8;bcd1<=2;bcd0<=2; end
			4823: begin bcd3<=4;bcd2<=8;bcd1<=2;bcd0<=3; end
			4824: begin bcd3<=4;bcd2<=8;bcd1<=2;bcd0<=4; end
			4825: begin bcd3<=4;bcd2<=8;bcd1<=2;bcd0<=5; end
			4826: begin bcd3<=4;bcd2<=8;bcd1<=2;bcd0<=6; end
			4827: begin bcd3<=4;bcd2<=8;bcd1<=2;bcd0<=7; end
			4828: begin bcd3<=4;bcd2<=8;bcd1<=2;bcd0<=8; end
			4829: begin bcd3<=4;bcd2<=8;bcd1<=2;bcd0<=9; end
			4830: begin bcd3<=4;bcd2<=8;bcd1<=3;bcd0<=0; end
			4831: begin bcd3<=4;bcd2<=8;bcd1<=3;bcd0<=1; end
			4832: begin bcd3<=4;bcd2<=8;bcd1<=3;bcd0<=2; end
			4833: begin bcd3<=4;bcd2<=8;bcd1<=3;bcd0<=3; end
			4834: begin bcd3<=4;bcd2<=8;bcd1<=3;bcd0<=4; end
			4835: begin bcd3<=4;bcd2<=8;bcd1<=3;bcd0<=5; end
			4836: begin bcd3<=4;bcd2<=8;bcd1<=3;bcd0<=6; end
			4837: begin bcd3<=4;bcd2<=8;bcd1<=3;bcd0<=7; end
			4838: begin bcd3<=4;bcd2<=8;bcd1<=3;bcd0<=8; end
			4839: begin bcd3<=4;bcd2<=8;bcd1<=3;bcd0<=9; end
			4840: begin bcd3<=4;bcd2<=8;bcd1<=4;bcd0<=0; end
			4841: begin bcd3<=4;bcd2<=8;bcd1<=4;bcd0<=1; end
			4842: begin bcd3<=4;bcd2<=8;bcd1<=4;bcd0<=2; end
			4843: begin bcd3<=4;bcd2<=8;bcd1<=4;bcd0<=3; end
			4844: begin bcd3<=4;bcd2<=8;bcd1<=4;bcd0<=4; end
			4845: begin bcd3<=4;bcd2<=8;bcd1<=4;bcd0<=5; end
			4846: begin bcd3<=4;bcd2<=8;bcd1<=4;bcd0<=6; end
			4847: begin bcd3<=4;bcd2<=8;bcd1<=4;bcd0<=7; end
			4848: begin bcd3<=4;bcd2<=8;bcd1<=4;bcd0<=8; end
			4849: begin bcd3<=4;bcd2<=8;bcd1<=4;bcd0<=9; end
			4850: begin bcd3<=4;bcd2<=8;bcd1<=5;bcd0<=0; end
			4851: begin bcd3<=4;bcd2<=8;bcd1<=5;bcd0<=1; end
			4852: begin bcd3<=4;bcd2<=8;bcd1<=5;bcd0<=2; end
			4853: begin bcd3<=4;bcd2<=8;bcd1<=5;bcd0<=3; end
			4854: begin bcd3<=4;bcd2<=8;bcd1<=5;bcd0<=4; end
			4855: begin bcd3<=4;bcd2<=8;bcd1<=5;bcd0<=5; end
			4856: begin bcd3<=4;bcd2<=8;bcd1<=5;bcd0<=6; end
			4857: begin bcd3<=4;bcd2<=8;bcd1<=5;bcd0<=7; end
			4858: begin bcd3<=4;bcd2<=8;bcd1<=5;bcd0<=8; end
			4859: begin bcd3<=4;bcd2<=8;bcd1<=5;bcd0<=9; end
			4860: begin bcd3<=4;bcd2<=8;bcd1<=6;bcd0<=0; end
			4861: begin bcd3<=4;bcd2<=8;bcd1<=6;bcd0<=1; end
			4862: begin bcd3<=4;bcd2<=8;bcd1<=6;bcd0<=2; end
			4863: begin bcd3<=4;bcd2<=8;bcd1<=6;bcd0<=3; end
			4864: begin bcd3<=4;bcd2<=8;bcd1<=6;bcd0<=4; end
			4865: begin bcd3<=4;bcd2<=8;bcd1<=6;bcd0<=5; end
			4866: begin bcd3<=4;bcd2<=8;bcd1<=6;bcd0<=6; end
			4867: begin bcd3<=4;bcd2<=8;bcd1<=6;bcd0<=7; end
			4868: begin bcd3<=4;bcd2<=8;bcd1<=6;bcd0<=8; end
			4869: begin bcd3<=4;bcd2<=8;bcd1<=6;bcd0<=9; end
			4870: begin bcd3<=4;bcd2<=8;bcd1<=7;bcd0<=0; end
			4871: begin bcd3<=4;bcd2<=8;bcd1<=7;bcd0<=1; end
			4872: begin bcd3<=4;bcd2<=8;bcd1<=7;bcd0<=2; end
			4873: begin bcd3<=4;bcd2<=8;bcd1<=7;bcd0<=3; end
			4874: begin bcd3<=4;bcd2<=8;bcd1<=7;bcd0<=4; end
			4875: begin bcd3<=4;bcd2<=8;bcd1<=7;bcd0<=5; end
			4876: begin bcd3<=4;bcd2<=8;bcd1<=7;bcd0<=6; end
			4877: begin bcd3<=4;bcd2<=8;bcd1<=7;bcd0<=7; end
			4878: begin bcd3<=4;bcd2<=8;bcd1<=7;bcd0<=8; end
			4879: begin bcd3<=4;bcd2<=8;bcd1<=7;bcd0<=9; end
			4880: begin bcd3<=4;bcd2<=8;bcd1<=8;bcd0<=0; end
			4881: begin bcd3<=4;bcd2<=8;bcd1<=8;bcd0<=1; end
			4882: begin bcd3<=4;bcd2<=8;bcd1<=8;bcd0<=2; end
			4883: begin bcd3<=4;bcd2<=8;bcd1<=8;bcd0<=3; end
			4884: begin bcd3<=4;bcd2<=8;bcd1<=8;bcd0<=4; end
			4885: begin bcd3<=4;bcd2<=8;bcd1<=8;bcd0<=5; end
			4886: begin bcd3<=4;bcd2<=8;bcd1<=8;bcd0<=6; end
			4887: begin bcd3<=4;bcd2<=8;bcd1<=8;bcd0<=7; end
			4888: begin bcd3<=4;bcd2<=8;bcd1<=8;bcd0<=8; end
			4889: begin bcd3<=4;bcd2<=8;bcd1<=8;bcd0<=9; end
			4890: begin bcd3<=4;bcd2<=8;bcd1<=9;bcd0<=0; end
			4891: begin bcd3<=4;bcd2<=8;bcd1<=9;bcd0<=1; end
			4892: begin bcd3<=4;bcd2<=8;bcd1<=9;bcd0<=2; end
			4893: begin bcd3<=4;bcd2<=8;bcd1<=9;bcd0<=3; end
			4894: begin bcd3<=4;bcd2<=8;bcd1<=9;bcd0<=4; end
			4895: begin bcd3<=4;bcd2<=8;bcd1<=9;bcd0<=5; end
			4896: begin bcd3<=4;bcd2<=8;bcd1<=9;bcd0<=6; end
			4897: begin bcd3<=4;bcd2<=8;bcd1<=9;bcd0<=7; end
			4898: begin bcd3<=4;bcd2<=8;bcd1<=9;bcd0<=8; end
			4899: begin bcd3<=4;bcd2<=8;bcd1<=9;bcd0<=9; end
			4900: begin bcd3<=4;bcd2<=9;bcd1<=0;bcd0<=0; end
			4901: begin bcd3<=4;bcd2<=9;bcd1<=0;bcd0<=1; end
			4902: begin bcd3<=4;bcd2<=9;bcd1<=0;bcd0<=2; end
			4903: begin bcd3<=4;bcd2<=9;bcd1<=0;bcd0<=3; end
			4904: begin bcd3<=4;bcd2<=9;bcd1<=0;bcd0<=4; end
			4905: begin bcd3<=4;bcd2<=9;bcd1<=0;bcd0<=5; end
			4906: begin bcd3<=4;bcd2<=9;bcd1<=0;bcd0<=6; end
			4907: begin bcd3<=4;bcd2<=9;bcd1<=0;bcd0<=7; end
			4908: begin bcd3<=4;bcd2<=9;bcd1<=0;bcd0<=8; end
			4909: begin bcd3<=4;bcd2<=9;bcd1<=0;bcd0<=9; end
			4910: begin bcd3<=4;bcd2<=9;bcd1<=1;bcd0<=0; end
			4911: begin bcd3<=4;bcd2<=9;bcd1<=1;bcd0<=1; end
			4912: begin bcd3<=4;bcd2<=9;bcd1<=1;bcd0<=2; end
			4913: begin bcd3<=4;bcd2<=9;bcd1<=1;bcd0<=3; end
			4914: begin bcd3<=4;bcd2<=9;bcd1<=1;bcd0<=4; end
			4915: begin bcd3<=4;bcd2<=9;bcd1<=1;bcd0<=5; end
			4916: begin bcd3<=4;bcd2<=9;bcd1<=1;bcd0<=6; end
			4917: begin bcd3<=4;bcd2<=9;bcd1<=1;bcd0<=7; end
			4918: begin bcd3<=4;bcd2<=9;bcd1<=1;bcd0<=8; end
			4919: begin bcd3<=4;bcd2<=9;bcd1<=1;bcd0<=9; end
			4920: begin bcd3<=4;bcd2<=9;bcd1<=2;bcd0<=0; end
			4921: begin bcd3<=4;bcd2<=9;bcd1<=2;bcd0<=1; end
			4922: begin bcd3<=4;bcd2<=9;bcd1<=2;bcd0<=2; end
			4923: begin bcd3<=4;bcd2<=9;bcd1<=2;bcd0<=3; end
			4924: begin bcd3<=4;bcd2<=9;bcd1<=2;bcd0<=4; end
			4925: begin bcd3<=4;bcd2<=9;bcd1<=2;bcd0<=5; end
			4926: begin bcd3<=4;bcd2<=9;bcd1<=2;bcd0<=6; end
			4927: begin bcd3<=4;bcd2<=9;bcd1<=2;bcd0<=7; end
			4928: begin bcd3<=4;bcd2<=9;bcd1<=2;bcd0<=8; end
			4929: begin bcd3<=4;bcd2<=9;bcd1<=2;bcd0<=9; end
			4930: begin bcd3<=4;bcd2<=9;bcd1<=3;bcd0<=0; end
			4931: begin bcd3<=4;bcd2<=9;bcd1<=3;bcd0<=1; end
			4932: begin bcd3<=4;bcd2<=9;bcd1<=3;bcd0<=2; end
			4933: begin bcd3<=4;bcd2<=9;bcd1<=3;bcd0<=3; end
			4934: begin bcd3<=4;bcd2<=9;bcd1<=3;bcd0<=4; end
			4935: begin bcd3<=4;bcd2<=9;bcd1<=3;bcd0<=5; end
			4936: begin bcd3<=4;bcd2<=9;bcd1<=3;bcd0<=6; end
			4937: begin bcd3<=4;bcd2<=9;bcd1<=3;bcd0<=7; end
			4938: begin bcd3<=4;bcd2<=9;bcd1<=3;bcd0<=8; end
			4939: begin bcd3<=4;bcd2<=9;bcd1<=3;bcd0<=9; end
			4940: begin bcd3<=4;bcd2<=9;bcd1<=4;bcd0<=0; end
			4941: begin bcd3<=4;bcd2<=9;bcd1<=4;bcd0<=1; end
			4942: begin bcd3<=4;bcd2<=9;bcd1<=4;bcd0<=2; end
			4943: begin bcd3<=4;bcd2<=9;bcd1<=4;bcd0<=3; end
			4944: begin bcd3<=4;bcd2<=9;bcd1<=4;bcd0<=4; end
			4945: begin bcd3<=4;bcd2<=9;bcd1<=4;bcd0<=5; end
			4946: begin bcd3<=4;bcd2<=9;bcd1<=4;bcd0<=6; end
			4947: begin bcd3<=4;bcd2<=9;bcd1<=4;bcd0<=7; end
			4948: begin bcd3<=4;bcd2<=9;bcd1<=4;bcd0<=8; end
			4949: begin bcd3<=4;bcd2<=9;bcd1<=4;bcd0<=9; end
			4950: begin bcd3<=4;bcd2<=9;bcd1<=5;bcd0<=0; end
			4951: begin bcd3<=4;bcd2<=9;bcd1<=5;bcd0<=1; end
			4952: begin bcd3<=4;bcd2<=9;bcd1<=5;bcd0<=2; end
			4953: begin bcd3<=4;bcd2<=9;bcd1<=5;bcd0<=3; end
			4954: begin bcd3<=4;bcd2<=9;bcd1<=5;bcd0<=4; end
			4955: begin bcd3<=4;bcd2<=9;bcd1<=5;bcd0<=5; end
			4956: begin bcd3<=4;bcd2<=9;bcd1<=5;bcd0<=6; end
			4957: begin bcd3<=4;bcd2<=9;bcd1<=5;bcd0<=7; end
			4958: begin bcd3<=4;bcd2<=9;bcd1<=5;bcd0<=8; end
			4959: begin bcd3<=4;bcd2<=9;bcd1<=5;bcd0<=9; end
			4960: begin bcd3<=4;bcd2<=9;bcd1<=6;bcd0<=0; end
			4961: begin bcd3<=4;bcd2<=9;bcd1<=6;bcd0<=1; end
			4962: begin bcd3<=4;bcd2<=9;bcd1<=6;bcd0<=2; end
			4963: begin bcd3<=4;bcd2<=9;bcd1<=6;bcd0<=3; end
			4964: begin bcd3<=4;bcd2<=9;bcd1<=6;bcd0<=4; end
			4965: begin bcd3<=4;bcd2<=9;bcd1<=6;bcd0<=5; end
			4966: begin bcd3<=4;bcd2<=9;bcd1<=6;bcd0<=6; end
			4967: begin bcd3<=4;bcd2<=9;bcd1<=6;bcd0<=7; end
			4968: begin bcd3<=4;bcd2<=9;bcd1<=6;bcd0<=8; end
			4969: begin bcd3<=4;bcd2<=9;bcd1<=6;bcd0<=9; end
			4970: begin bcd3<=4;bcd2<=9;bcd1<=7;bcd0<=0; end
			4971: begin bcd3<=4;bcd2<=9;bcd1<=7;bcd0<=1; end
			4972: begin bcd3<=4;bcd2<=9;bcd1<=7;bcd0<=2; end
			4973: begin bcd3<=4;bcd2<=9;bcd1<=7;bcd0<=3; end
			4974: begin bcd3<=4;bcd2<=9;bcd1<=7;bcd0<=4; end
			4975: begin bcd3<=4;bcd2<=9;bcd1<=7;bcd0<=5; end
			4976: begin bcd3<=4;bcd2<=9;bcd1<=7;bcd0<=6; end
			4977: begin bcd3<=4;bcd2<=9;bcd1<=7;bcd0<=7; end
			4978: begin bcd3<=4;bcd2<=9;bcd1<=7;bcd0<=8; end
			4979: begin bcd3<=4;bcd2<=9;bcd1<=7;bcd0<=9; end
			4980: begin bcd3<=4;bcd2<=9;bcd1<=8;bcd0<=0; end
			4981: begin bcd3<=4;bcd2<=9;bcd1<=8;bcd0<=1; end
			4982: begin bcd3<=4;bcd2<=9;bcd1<=8;bcd0<=2; end
			4983: begin bcd3<=4;bcd2<=9;bcd1<=8;bcd0<=3; end
			4984: begin bcd3<=4;bcd2<=9;bcd1<=8;bcd0<=4; end
			4985: begin bcd3<=4;bcd2<=9;bcd1<=8;bcd0<=5; end
			4986: begin bcd3<=4;bcd2<=9;bcd1<=8;bcd0<=6; end
			4987: begin bcd3<=4;bcd2<=9;bcd1<=8;bcd0<=7; end
			4988: begin bcd3<=4;bcd2<=9;bcd1<=8;bcd0<=8; end
			4989: begin bcd3<=4;bcd2<=9;bcd1<=8;bcd0<=9; end
			4990: begin bcd3<=4;bcd2<=9;bcd1<=9;bcd0<=0; end
			4991: begin bcd3<=4;bcd2<=9;bcd1<=9;bcd0<=1; end
			4992: begin bcd3<=4;bcd2<=9;bcd1<=9;bcd0<=2; end
			4993: begin bcd3<=4;bcd2<=9;bcd1<=9;bcd0<=3; end
			4994: begin bcd3<=4;bcd2<=9;bcd1<=9;bcd0<=4; end
			4995: begin bcd3<=4;bcd2<=9;bcd1<=9;bcd0<=5; end
			4996: begin bcd3<=4;bcd2<=9;bcd1<=9;bcd0<=6; end
			4997: begin bcd3<=4;bcd2<=9;bcd1<=9;bcd0<=7; end
			4998: begin bcd3<=4;bcd2<=9;bcd1<=9;bcd0<=8; end
			4999: begin bcd3<=4;bcd2<=9;bcd1<=9;bcd0<=9; end
			5000: begin bcd3<=5;bcd2<=0;bcd1<=0;bcd0<=0; end
			5001: begin bcd3<=5;bcd2<=0;bcd1<=0;bcd0<=1; end
			5002: begin bcd3<=5;bcd2<=0;bcd1<=0;bcd0<=2; end
			5003: begin bcd3<=5;bcd2<=0;bcd1<=0;bcd0<=3; end
			5004: begin bcd3<=5;bcd2<=0;bcd1<=0;bcd0<=4; end
			5005: begin bcd3<=5;bcd2<=0;bcd1<=0;bcd0<=5; end
			5006: begin bcd3<=5;bcd2<=0;bcd1<=0;bcd0<=6; end
			5007: begin bcd3<=5;bcd2<=0;bcd1<=0;bcd0<=7; end
			5008: begin bcd3<=5;bcd2<=0;bcd1<=0;bcd0<=8; end
			5009: begin bcd3<=5;bcd2<=0;bcd1<=0;bcd0<=9; end
			5010: begin bcd3<=5;bcd2<=0;bcd1<=1;bcd0<=0; end
			5011: begin bcd3<=5;bcd2<=0;bcd1<=1;bcd0<=1; end
			5012: begin bcd3<=5;bcd2<=0;bcd1<=1;bcd0<=2; end
			5013: begin bcd3<=5;bcd2<=0;bcd1<=1;bcd0<=3; end
			5014: begin bcd3<=5;bcd2<=0;bcd1<=1;bcd0<=4; end
			5015: begin bcd3<=5;bcd2<=0;bcd1<=1;bcd0<=5; end
			5016: begin bcd3<=5;bcd2<=0;bcd1<=1;bcd0<=6; end
			5017: begin bcd3<=5;bcd2<=0;bcd1<=1;bcd0<=7; end
			5018: begin bcd3<=5;bcd2<=0;bcd1<=1;bcd0<=8; end
			5019: begin bcd3<=5;bcd2<=0;bcd1<=1;bcd0<=9; end
			5020: begin bcd3<=5;bcd2<=0;bcd1<=2;bcd0<=0; end
			5021: begin bcd3<=5;bcd2<=0;bcd1<=2;bcd0<=1; end
			5022: begin bcd3<=5;bcd2<=0;bcd1<=2;bcd0<=2; end
			5023: begin bcd3<=5;bcd2<=0;bcd1<=2;bcd0<=3; end
			5024: begin bcd3<=5;bcd2<=0;bcd1<=2;bcd0<=4; end
			5025: begin bcd3<=5;bcd2<=0;bcd1<=2;bcd0<=5; end
			5026: begin bcd3<=5;bcd2<=0;bcd1<=2;bcd0<=6; end
			5027: begin bcd3<=5;bcd2<=0;bcd1<=2;bcd0<=7; end
			5028: begin bcd3<=5;bcd2<=0;bcd1<=2;bcd0<=8; end
			5029: begin bcd3<=5;bcd2<=0;bcd1<=2;bcd0<=9; end
			5030: begin bcd3<=5;bcd2<=0;bcd1<=3;bcd0<=0; end
			5031: begin bcd3<=5;bcd2<=0;bcd1<=3;bcd0<=1; end
			5032: begin bcd3<=5;bcd2<=0;bcd1<=3;bcd0<=2; end
			5033: begin bcd3<=5;bcd2<=0;bcd1<=3;bcd0<=3; end
			5034: begin bcd3<=5;bcd2<=0;bcd1<=3;bcd0<=4; end
			5035: begin bcd3<=5;bcd2<=0;bcd1<=3;bcd0<=5; end
			5036: begin bcd3<=5;bcd2<=0;bcd1<=3;bcd0<=6; end
			5037: begin bcd3<=5;bcd2<=0;bcd1<=3;bcd0<=7; end
			5038: begin bcd3<=5;bcd2<=0;bcd1<=3;bcd0<=8; end
			5039: begin bcd3<=5;bcd2<=0;bcd1<=3;bcd0<=9; end
			5040: begin bcd3<=5;bcd2<=0;bcd1<=4;bcd0<=0; end
			5041: begin bcd3<=5;bcd2<=0;bcd1<=4;bcd0<=1; end
			5042: begin bcd3<=5;bcd2<=0;bcd1<=4;bcd0<=2; end
			5043: begin bcd3<=5;bcd2<=0;bcd1<=4;bcd0<=3; end
			5044: begin bcd3<=5;bcd2<=0;bcd1<=4;bcd0<=4; end
			5045: begin bcd3<=5;bcd2<=0;bcd1<=4;bcd0<=5; end
			5046: begin bcd3<=5;bcd2<=0;bcd1<=4;bcd0<=6; end
			5047: begin bcd3<=5;bcd2<=0;bcd1<=4;bcd0<=7; end
			5048: begin bcd3<=5;bcd2<=0;bcd1<=4;bcd0<=8; end
			5049: begin bcd3<=5;bcd2<=0;bcd1<=4;bcd0<=9; end
			5050: begin bcd3<=5;bcd2<=0;bcd1<=5;bcd0<=0; end
			5051: begin bcd3<=5;bcd2<=0;bcd1<=5;bcd0<=1; end
			5052: begin bcd3<=5;bcd2<=0;bcd1<=5;bcd0<=2; end
			5053: begin bcd3<=5;bcd2<=0;bcd1<=5;bcd0<=3; end
			5054: begin bcd3<=5;bcd2<=0;bcd1<=5;bcd0<=4; end
			5055: begin bcd3<=5;bcd2<=0;bcd1<=5;bcd0<=5; end
			5056: begin bcd3<=5;bcd2<=0;bcd1<=5;bcd0<=6; end
			5057: begin bcd3<=5;bcd2<=0;bcd1<=5;bcd0<=7; end
			5058: begin bcd3<=5;bcd2<=0;bcd1<=5;bcd0<=8; end
			5059: begin bcd3<=5;bcd2<=0;bcd1<=5;bcd0<=9; end
			5060: begin bcd3<=5;bcd2<=0;bcd1<=6;bcd0<=0; end
			5061: begin bcd3<=5;bcd2<=0;bcd1<=6;bcd0<=1; end
			5062: begin bcd3<=5;bcd2<=0;bcd1<=6;bcd0<=2; end
			5063: begin bcd3<=5;bcd2<=0;bcd1<=6;bcd0<=3; end
			5064: begin bcd3<=5;bcd2<=0;bcd1<=6;bcd0<=4; end
			5065: begin bcd3<=5;bcd2<=0;bcd1<=6;bcd0<=5; end
			5066: begin bcd3<=5;bcd2<=0;bcd1<=6;bcd0<=6; end
			5067: begin bcd3<=5;bcd2<=0;bcd1<=6;bcd0<=7; end
			5068: begin bcd3<=5;bcd2<=0;bcd1<=6;bcd0<=8; end
			5069: begin bcd3<=5;bcd2<=0;bcd1<=6;bcd0<=9; end
			5070: begin bcd3<=5;bcd2<=0;bcd1<=7;bcd0<=0; end
			5071: begin bcd3<=5;bcd2<=0;bcd1<=7;bcd0<=1; end
			5072: begin bcd3<=5;bcd2<=0;bcd1<=7;bcd0<=2; end
			5073: begin bcd3<=5;bcd2<=0;bcd1<=7;bcd0<=3; end
			5074: begin bcd3<=5;bcd2<=0;bcd1<=7;bcd0<=4; end
			5075: begin bcd3<=5;bcd2<=0;bcd1<=7;bcd0<=5; end
			5076: begin bcd3<=5;bcd2<=0;bcd1<=7;bcd0<=6; end
			5077: begin bcd3<=5;bcd2<=0;bcd1<=7;bcd0<=7; end
			5078: begin bcd3<=5;bcd2<=0;bcd1<=7;bcd0<=8; end
			5079: begin bcd3<=5;bcd2<=0;bcd1<=7;bcd0<=9; end
			5080: begin bcd3<=5;bcd2<=0;bcd1<=8;bcd0<=0; end
			5081: begin bcd3<=5;bcd2<=0;bcd1<=8;bcd0<=1; end
			5082: begin bcd3<=5;bcd2<=0;bcd1<=8;bcd0<=2; end
			5083: begin bcd3<=5;bcd2<=0;bcd1<=8;bcd0<=3; end
			5084: begin bcd3<=5;bcd2<=0;bcd1<=8;bcd0<=4; end
			5085: begin bcd3<=5;bcd2<=0;bcd1<=8;bcd0<=5; end
			5086: begin bcd3<=5;bcd2<=0;bcd1<=8;bcd0<=6; end
			5087: begin bcd3<=5;bcd2<=0;bcd1<=8;bcd0<=7; end
			5088: begin bcd3<=5;bcd2<=0;bcd1<=8;bcd0<=8; end
			5089: begin bcd3<=5;bcd2<=0;bcd1<=8;bcd0<=9; end
			5090: begin bcd3<=5;bcd2<=0;bcd1<=9;bcd0<=0; end
			5091: begin bcd3<=5;bcd2<=0;bcd1<=9;bcd0<=1; end
			5092: begin bcd3<=5;bcd2<=0;bcd1<=9;bcd0<=2; end
			5093: begin bcd3<=5;bcd2<=0;bcd1<=9;bcd0<=3; end
			5094: begin bcd3<=5;bcd2<=0;bcd1<=9;bcd0<=4; end
			5095: begin bcd3<=5;bcd2<=0;bcd1<=9;bcd0<=5; end
			5096: begin bcd3<=5;bcd2<=0;bcd1<=9;bcd0<=6; end
			5097: begin bcd3<=5;bcd2<=0;bcd1<=9;bcd0<=7; end
			5098: begin bcd3<=5;bcd2<=0;bcd1<=9;bcd0<=8; end
			5099: begin bcd3<=5;bcd2<=0;bcd1<=9;bcd0<=9; end
			5100: begin bcd3<=5;bcd2<=1;bcd1<=0;bcd0<=0; end
			5101: begin bcd3<=5;bcd2<=1;bcd1<=0;bcd0<=1; end
			5102: begin bcd3<=5;bcd2<=1;bcd1<=0;bcd0<=2; end
			5103: begin bcd3<=5;bcd2<=1;bcd1<=0;bcd0<=3; end
			5104: begin bcd3<=5;bcd2<=1;bcd1<=0;bcd0<=4; end
			5105: begin bcd3<=5;bcd2<=1;bcd1<=0;bcd0<=5; end
			5106: begin bcd3<=5;bcd2<=1;bcd1<=0;bcd0<=6; end
			5107: begin bcd3<=5;bcd2<=1;bcd1<=0;bcd0<=7; end
			5108: begin bcd3<=5;bcd2<=1;bcd1<=0;bcd0<=8; end
			5109: begin bcd3<=5;bcd2<=1;bcd1<=0;bcd0<=9; end
			5110: begin bcd3<=5;bcd2<=1;bcd1<=1;bcd0<=0; end
			5111: begin bcd3<=5;bcd2<=1;bcd1<=1;bcd0<=1; end
			5112: begin bcd3<=5;bcd2<=1;bcd1<=1;bcd0<=2; end
			5113: begin bcd3<=5;bcd2<=1;bcd1<=1;bcd0<=3; end
			5114: begin bcd3<=5;bcd2<=1;bcd1<=1;bcd0<=4; end
			5115: begin bcd3<=5;bcd2<=1;bcd1<=1;bcd0<=5; end
			5116: begin bcd3<=5;bcd2<=1;bcd1<=1;bcd0<=6; end
			5117: begin bcd3<=5;bcd2<=1;bcd1<=1;bcd0<=7; end
			5118: begin bcd3<=5;bcd2<=1;bcd1<=1;bcd0<=8; end
			5119: begin bcd3<=5;bcd2<=1;bcd1<=1;bcd0<=9; end
			5120: begin bcd3<=5;bcd2<=1;bcd1<=2;bcd0<=0; end
			5121: begin bcd3<=5;bcd2<=1;bcd1<=2;bcd0<=1; end
			5122: begin bcd3<=5;bcd2<=1;bcd1<=2;bcd0<=2; end
			5123: begin bcd3<=5;bcd2<=1;bcd1<=2;bcd0<=3; end
			5124: begin bcd3<=5;bcd2<=1;bcd1<=2;bcd0<=4; end
			5125: begin bcd3<=5;bcd2<=1;bcd1<=2;bcd0<=5; end
			5126: begin bcd3<=5;bcd2<=1;bcd1<=2;bcd0<=6; end
			5127: begin bcd3<=5;bcd2<=1;bcd1<=2;bcd0<=7; end
			5128: begin bcd3<=5;bcd2<=1;bcd1<=2;bcd0<=8; end
			5129: begin bcd3<=5;bcd2<=1;bcd1<=2;bcd0<=9; end
			5130: begin bcd3<=5;bcd2<=1;bcd1<=3;bcd0<=0; end
			5131: begin bcd3<=5;bcd2<=1;bcd1<=3;bcd0<=1; end
			5132: begin bcd3<=5;bcd2<=1;bcd1<=3;bcd0<=2; end
			5133: begin bcd3<=5;bcd2<=1;bcd1<=3;bcd0<=3; end
			5134: begin bcd3<=5;bcd2<=1;bcd1<=3;bcd0<=4; end
			5135: begin bcd3<=5;bcd2<=1;bcd1<=3;bcd0<=5; end
			5136: begin bcd3<=5;bcd2<=1;bcd1<=3;bcd0<=6; end
			5137: begin bcd3<=5;bcd2<=1;bcd1<=3;bcd0<=7; end
			5138: begin bcd3<=5;bcd2<=1;bcd1<=3;bcd0<=8; end
			5139: begin bcd3<=5;bcd2<=1;bcd1<=3;bcd0<=9; end
			5140: begin bcd3<=5;bcd2<=1;bcd1<=4;bcd0<=0; end
			5141: begin bcd3<=5;bcd2<=1;bcd1<=4;bcd0<=1; end
			5142: begin bcd3<=5;bcd2<=1;bcd1<=4;bcd0<=2; end
			5143: begin bcd3<=5;bcd2<=1;bcd1<=4;bcd0<=3; end
			5144: begin bcd3<=5;bcd2<=1;bcd1<=4;bcd0<=4; end
			5145: begin bcd3<=5;bcd2<=1;bcd1<=4;bcd0<=5; end
			5146: begin bcd3<=5;bcd2<=1;bcd1<=4;bcd0<=6; end
			5147: begin bcd3<=5;bcd2<=1;bcd1<=4;bcd0<=7; end
			5148: begin bcd3<=5;bcd2<=1;bcd1<=4;bcd0<=8; end
			5149: begin bcd3<=5;bcd2<=1;bcd1<=4;bcd0<=9; end
			5150: begin bcd3<=5;bcd2<=1;bcd1<=5;bcd0<=0; end
			5151: begin bcd3<=5;bcd2<=1;bcd1<=5;bcd0<=1; end
			5152: begin bcd3<=5;bcd2<=1;bcd1<=5;bcd0<=2; end
			5153: begin bcd3<=5;bcd2<=1;bcd1<=5;bcd0<=3; end
			5154: begin bcd3<=5;bcd2<=1;bcd1<=5;bcd0<=4; end
			5155: begin bcd3<=5;bcd2<=1;bcd1<=5;bcd0<=5; end
			5156: begin bcd3<=5;bcd2<=1;bcd1<=5;bcd0<=6; end
			5157: begin bcd3<=5;bcd2<=1;bcd1<=5;bcd0<=7; end
			5158: begin bcd3<=5;bcd2<=1;bcd1<=5;bcd0<=8; end
			5159: begin bcd3<=5;bcd2<=1;bcd1<=5;bcd0<=9; end
			5160: begin bcd3<=5;bcd2<=1;bcd1<=6;bcd0<=0; end
			5161: begin bcd3<=5;bcd2<=1;bcd1<=6;bcd0<=1; end
			5162: begin bcd3<=5;bcd2<=1;bcd1<=6;bcd0<=2; end
			5163: begin bcd3<=5;bcd2<=1;bcd1<=6;bcd0<=3; end
			5164: begin bcd3<=5;bcd2<=1;bcd1<=6;bcd0<=4; end
			5165: begin bcd3<=5;bcd2<=1;bcd1<=6;bcd0<=5; end
			5166: begin bcd3<=5;bcd2<=1;bcd1<=6;bcd0<=6; end
			5167: begin bcd3<=5;bcd2<=1;bcd1<=6;bcd0<=7; end
			5168: begin bcd3<=5;bcd2<=1;bcd1<=6;bcd0<=8; end
			5169: begin bcd3<=5;bcd2<=1;bcd1<=6;bcd0<=9; end
			5170: begin bcd3<=5;bcd2<=1;bcd1<=7;bcd0<=0; end
			5171: begin bcd3<=5;bcd2<=1;bcd1<=7;bcd0<=1; end
			5172: begin bcd3<=5;bcd2<=1;bcd1<=7;bcd0<=2; end
			5173: begin bcd3<=5;bcd2<=1;bcd1<=7;bcd0<=3; end
			5174: begin bcd3<=5;bcd2<=1;bcd1<=7;bcd0<=4; end
			5175: begin bcd3<=5;bcd2<=1;bcd1<=7;bcd0<=5; end
			5176: begin bcd3<=5;bcd2<=1;bcd1<=7;bcd0<=6; end
			5177: begin bcd3<=5;bcd2<=1;bcd1<=7;bcd0<=7; end
			5178: begin bcd3<=5;bcd2<=1;bcd1<=7;bcd0<=8; end
			5179: begin bcd3<=5;bcd2<=1;bcd1<=7;bcd0<=9; end
			5180: begin bcd3<=5;bcd2<=1;bcd1<=8;bcd0<=0; end
			5181: begin bcd3<=5;bcd2<=1;bcd1<=8;bcd0<=1; end
			5182: begin bcd3<=5;bcd2<=1;bcd1<=8;bcd0<=2; end
			5183: begin bcd3<=5;bcd2<=1;bcd1<=8;bcd0<=3; end
			5184: begin bcd3<=5;bcd2<=1;bcd1<=8;bcd0<=4; end
			5185: begin bcd3<=5;bcd2<=1;bcd1<=8;bcd0<=5; end
			5186: begin bcd3<=5;bcd2<=1;bcd1<=8;bcd0<=6; end
			5187: begin bcd3<=5;bcd2<=1;bcd1<=8;bcd0<=7; end
			5188: begin bcd3<=5;bcd2<=1;bcd1<=8;bcd0<=8; end
			5189: begin bcd3<=5;bcd2<=1;bcd1<=8;bcd0<=9; end
			5190: begin bcd3<=5;bcd2<=1;bcd1<=9;bcd0<=0; end
			5191: begin bcd3<=5;bcd2<=1;bcd1<=9;bcd0<=1; end
			5192: begin bcd3<=5;bcd2<=1;bcd1<=9;bcd0<=2; end
			5193: begin bcd3<=5;bcd2<=1;bcd1<=9;bcd0<=3; end
			5194: begin bcd3<=5;bcd2<=1;bcd1<=9;bcd0<=4; end
			5195: begin bcd3<=5;bcd2<=1;bcd1<=9;bcd0<=5; end
			5196: begin bcd3<=5;bcd2<=1;bcd1<=9;bcd0<=6; end
			5197: begin bcd3<=5;bcd2<=1;bcd1<=9;bcd0<=7; end
			5198: begin bcd3<=5;bcd2<=1;bcd1<=9;bcd0<=8; end
			5199: begin bcd3<=5;bcd2<=1;bcd1<=9;bcd0<=9; end
			5200: begin bcd3<=5;bcd2<=2;bcd1<=0;bcd0<=0; end
			5201: begin bcd3<=5;bcd2<=2;bcd1<=0;bcd0<=1; end
			5202: begin bcd3<=5;bcd2<=2;bcd1<=0;bcd0<=2; end
			5203: begin bcd3<=5;bcd2<=2;bcd1<=0;bcd0<=3; end
			5204: begin bcd3<=5;bcd2<=2;bcd1<=0;bcd0<=4; end
			5205: begin bcd3<=5;bcd2<=2;bcd1<=0;bcd0<=5; end
			5206: begin bcd3<=5;bcd2<=2;bcd1<=0;bcd0<=6; end
			5207: begin bcd3<=5;bcd2<=2;bcd1<=0;bcd0<=7; end
			5208: begin bcd3<=5;bcd2<=2;bcd1<=0;bcd0<=8; end
			5209: begin bcd3<=5;bcd2<=2;bcd1<=0;bcd0<=9; end
			5210: begin bcd3<=5;bcd2<=2;bcd1<=1;bcd0<=0; end
			5211: begin bcd3<=5;bcd2<=2;bcd1<=1;bcd0<=1; end
			5212: begin bcd3<=5;bcd2<=2;bcd1<=1;bcd0<=2; end
			5213: begin bcd3<=5;bcd2<=2;bcd1<=1;bcd0<=3; end
			5214: begin bcd3<=5;bcd2<=2;bcd1<=1;bcd0<=4; end
			5215: begin bcd3<=5;bcd2<=2;bcd1<=1;bcd0<=5; end
			5216: begin bcd3<=5;bcd2<=2;bcd1<=1;bcd0<=6; end
			5217: begin bcd3<=5;bcd2<=2;bcd1<=1;bcd0<=7; end
			5218: begin bcd3<=5;bcd2<=2;bcd1<=1;bcd0<=8; end
			5219: begin bcd3<=5;bcd2<=2;bcd1<=1;bcd0<=9; end
			5220: begin bcd3<=5;bcd2<=2;bcd1<=2;bcd0<=0; end
			5221: begin bcd3<=5;bcd2<=2;bcd1<=2;bcd0<=1; end
			5222: begin bcd3<=5;bcd2<=2;bcd1<=2;bcd0<=2; end
			5223: begin bcd3<=5;bcd2<=2;bcd1<=2;bcd0<=3; end
			5224: begin bcd3<=5;bcd2<=2;bcd1<=2;bcd0<=4; end
			5225: begin bcd3<=5;bcd2<=2;bcd1<=2;bcd0<=5; end
			5226: begin bcd3<=5;bcd2<=2;bcd1<=2;bcd0<=6; end
			5227: begin bcd3<=5;bcd2<=2;bcd1<=2;bcd0<=7; end
			5228: begin bcd3<=5;bcd2<=2;bcd1<=2;bcd0<=8; end
			5229: begin bcd3<=5;bcd2<=2;bcd1<=2;bcd0<=9; end
			5230: begin bcd3<=5;bcd2<=2;bcd1<=3;bcd0<=0; end
			5231: begin bcd3<=5;bcd2<=2;bcd1<=3;bcd0<=1; end
			5232: begin bcd3<=5;bcd2<=2;bcd1<=3;bcd0<=2; end
			5233: begin bcd3<=5;bcd2<=2;bcd1<=3;bcd0<=3; end
			5234: begin bcd3<=5;bcd2<=2;bcd1<=3;bcd0<=4; end
			5235: begin bcd3<=5;bcd2<=2;bcd1<=3;bcd0<=5; end
			5236: begin bcd3<=5;bcd2<=2;bcd1<=3;bcd0<=6; end
			5237: begin bcd3<=5;bcd2<=2;bcd1<=3;bcd0<=7; end
			5238: begin bcd3<=5;bcd2<=2;bcd1<=3;bcd0<=8; end
			5239: begin bcd3<=5;bcd2<=2;bcd1<=3;bcd0<=9; end
			5240: begin bcd3<=5;bcd2<=2;bcd1<=4;bcd0<=0; end
			5241: begin bcd3<=5;bcd2<=2;bcd1<=4;bcd0<=1; end
			5242: begin bcd3<=5;bcd2<=2;bcd1<=4;bcd0<=2; end
			5243: begin bcd3<=5;bcd2<=2;bcd1<=4;bcd0<=3; end
			5244: begin bcd3<=5;bcd2<=2;bcd1<=4;bcd0<=4; end
			5245: begin bcd3<=5;bcd2<=2;bcd1<=4;bcd0<=5; end
			5246: begin bcd3<=5;bcd2<=2;bcd1<=4;bcd0<=6; end
			5247: begin bcd3<=5;bcd2<=2;bcd1<=4;bcd0<=7; end
			5248: begin bcd3<=5;bcd2<=2;bcd1<=4;bcd0<=8; end
			5249: begin bcd3<=5;bcd2<=2;bcd1<=4;bcd0<=9; end
			5250: begin bcd3<=5;bcd2<=2;bcd1<=5;bcd0<=0; end
			5251: begin bcd3<=5;bcd2<=2;bcd1<=5;bcd0<=1; end
			5252: begin bcd3<=5;bcd2<=2;bcd1<=5;bcd0<=2; end
			5253: begin bcd3<=5;bcd2<=2;bcd1<=5;bcd0<=3; end
			5254: begin bcd3<=5;bcd2<=2;bcd1<=5;bcd0<=4; end
			5255: begin bcd3<=5;bcd2<=2;bcd1<=5;bcd0<=5; end
			5256: begin bcd3<=5;bcd2<=2;bcd1<=5;bcd0<=6; end
			5257: begin bcd3<=5;bcd2<=2;bcd1<=5;bcd0<=7; end
			5258: begin bcd3<=5;bcd2<=2;bcd1<=5;bcd0<=8; end
			5259: begin bcd3<=5;bcd2<=2;bcd1<=5;bcd0<=9; end
			5260: begin bcd3<=5;bcd2<=2;bcd1<=6;bcd0<=0; end
			5261: begin bcd3<=5;bcd2<=2;bcd1<=6;bcd0<=1; end
			5262: begin bcd3<=5;bcd2<=2;bcd1<=6;bcd0<=2; end
			5263: begin bcd3<=5;bcd2<=2;bcd1<=6;bcd0<=3; end
			5264: begin bcd3<=5;bcd2<=2;bcd1<=6;bcd0<=4; end
			5265: begin bcd3<=5;bcd2<=2;bcd1<=6;bcd0<=5; end
			5266: begin bcd3<=5;bcd2<=2;bcd1<=6;bcd0<=6; end
			5267: begin bcd3<=5;bcd2<=2;bcd1<=6;bcd0<=7; end
			5268: begin bcd3<=5;bcd2<=2;bcd1<=6;bcd0<=8; end
			5269: begin bcd3<=5;bcd2<=2;bcd1<=6;bcd0<=9; end
			5270: begin bcd3<=5;bcd2<=2;bcd1<=7;bcd0<=0; end
			5271: begin bcd3<=5;bcd2<=2;bcd1<=7;bcd0<=1; end
			5272: begin bcd3<=5;bcd2<=2;bcd1<=7;bcd0<=2; end
			5273: begin bcd3<=5;bcd2<=2;bcd1<=7;bcd0<=3; end
			5274: begin bcd3<=5;bcd2<=2;bcd1<=7;bcd0<=4; end
			5275: begin bcd3<=5;bcd2<=2;bcd1<=7;bcd0<=5; end
			5276: begin bcd3<=5;bcd2<=2;bcd1<=7;bcd0<=6; end
			5277: begin bcd3<=5;bcd2<=2;bcd1<=7;bcd0<=7; end
			5278: begin bcd3<=5;bcd2<=2;bcd1<=7;bcd0<=8; end
			5279: begin bcd3<=5;bcd2<=2;bcd1<=7;bcd0<=9; end
			5280: begin bcd3<=5;bcd2<=2;bcd1<=8;bcd0<=0; end
			5281: begin bcd3<=5;bcd2<=2;bcd1<=8;bcd0<=1; end
			5282: begin bcd3<=5;bcd2<=2;bcd1<=8;bcd0<=2; end
			5283: begin bcd3<=5;bcd2<=2;bcd1<=8;bcd0<=3; end
			5284: begin bcd3<=5;bcd2<=2;bcd1<=8;bcd0<=4; end
			5285: begin bcd3<=5;bcd2<=2;bcd1<=8;bcd0<=5; end
			5286: begin bcd3<=5;bcd2<=2;bcd1<=8;bcd0<=6; end
			5287: begin bcd3<=5;bcd2<=2;bcd1<=8;bcd0<=7; end
			5288: begin bcd3<=5;bcd2<=2;bcd1<=8;bcd0<=8; end
			5289: begin bcd3<=5;bcd2<=2;bcd1<=8;bcd0<=9; end
			5290: begin bcd3<=5;bcd2<=2;bcd1<=9;bcd0<=0; end
			5291: begin bcd3<=5;bcd2<=2;bcd1<=9;bcd0<=1; end
			5292: begin bcd3<=5;bcd2<=2;bcd1<=9;bcd0<=2; end
			5293: begin bcd3<=5;bcd2<=2;bcd1<=9;bcd0<=3; end
			5294: begin bcd3<=5;bcd2<=2;bcd1<=9;bcd0<=4; end
			5295: begin bcd3<=5;bcd2<=2;bcd1<=9;bcd0<=5; end
			5296: begin bcd3<=5;bcd2<=2;bcd1<=9;bcd0<=6; end
			5297: begin bcd3<=5;bcd2<=2;bcd1<=9;bcd0<=7; end
			5298: begin bcd3<=5;bcd2<=2;bcd1<=9;bcd0<=8; end
			5299: begin bcd3<=5;bcd2<=2;bcd1<=9;bcd0<=9; end
			5300: begin bcd3<=5;bcd2<=3;bcd1<=0;bcd0<=0; end
			5301: begin bcd3<=5;bcd2<=3;bcd1<=0;bcd0<=1; end
			5302: begin bcd3<=5;bcd2<=3;bcd1<=0;bcd0<=2; end
			5303: begin bcd3<=5;bcd2<=3;bcd1<=0;bcd0<=3; end
			5304: begin bcd3<=5;bcd2<=3;bcd1<=0;bcd0<=4; end
			5305: begin bcd3<=5;bcd2<=3;bcd1<=0;bcd0<=5; end
			5306: begin bcd3<=5;bcd2<=3;bcd1<=0;bcd0<=6; end
			5307: begin bcd3<=5;bcd2<=3;bcd1<=0;bcd0<=7; end
			5308: begin bcd3<=5;bcd2<=3;bcd1<=0;bcd0<=8; end
			5309: begin bcd3<=5;bcd2<=3;bcd1<=0;bcd0<=9; end
			5310: begin bcd3<=5;bcd2<=3;bcd1<=1;bcd0<=0; end
			5311: begin bcd3<=5;bcd2<=3;bcd1<=1;bcd0<=1; end
			5312: begin bcd3<=5;bcd2<=3;bcd1<=1;bcd0<=2; end
			5313: begin bcd3<=5;bcd2<=3;bcd1<=1;bcd0<=3; end
			5314: begin bcd3<=5;bcd2<=3;bcd1<=1;bcd0<=4; end
			5315: begin bcd3<=5;bcd2<=3;bcd1<=1;bcd0<=5; end
			5316: begin bcd3<=5;bcd2<=3;bcd1<=1;bcd0<=6; end
			5317: begin bcd3<=5;bcd2<=3;bcd1<=1;bcd0<=7; end
			5318: begin bcd3<=5;bcd2<=3;bcd1<=1;bcd0<=8; end
			5319: begin bcd3<=5;bcd2<=3;bcd1<=1;bcd0<=9; end
			5320: begin bcd3<=5;bcd2<=3;bcd1<=2;bcd0<=0; end
			5321: begin bcd3<=5;bcd2<=3;bcd1<=2;bcd0<=1; end
			5322: begin bcd3<=5;bcd2<=3;bcd1<=2;bcd0<=2; end
			5323: begin bcd3<=5;bcd2<=3;bcd1<=2;bcd0<=3; end
			5324: begin bcd3<=5;bcd2<=3;bcd1<=2;bcd0<=4; end
			5325: begin bcd3<=5;bcd2<=3;bcd1<=2;bcd0<=5; end
			5326: begin bcd3<=5;bcd2<=3;bcd1<=2;bcd0<=6; end
			5327: begin bcd3<=5;bcd2<=3;bcd1<=2;bcd0<=7; end
			5328: begin bcd3<=5;bcd2<=3;bcd1<=2;bcd0<=8; end
			5329: begin bcd3<=5;bcd2<=3;bcd1<=2;bcd0<=9; end
			5330: begin bcd3<=5;bcd2<=3;bcd1<=3;bcd0<=0; end
			5331: begin bcd3<=5;bcd2<=3;bcd1<=3;bcd0<=1; end
			5332: begin bcd3<=5;bcd2<=3;bcd1<=3;bcd0<=2; end
			5333: begin bcd3<=5;bcd2<=3;bcd1<=3;bcd0<=3; end
			5334: begin bcd3<=5;bcd2<=3;bcd1<=3;bcd0<=4; end
			5335: begin bcd3<=5;bcd2<=3;bcd1<=3;bcd0<=5; end
			5336: begin bcd3<=5;bcd2<=3;bcd1<=3;bcd0<=6; end
			5337: begin bcd3<=5;bcd2<=3;bcd1<=3;bcd0<=7; end
			5338: begin bcd3<=5;bcd2<=3;bcd1<=3;bcd0<=8; end
			5339: begin bcd3<=5;bcd2<=3;bcd1<=3;bcd0<=9; end
			5340: begin bcd3<=5;bcd2<=3;bcd1<=4;bcd0<=0; end
			5341: begin bcd3<=5;bcd2<=3;bcd1<=4;bcd0<=1; end
			5342: begin bcd3<=5;bcd2<=3;bcd1<=4;bcd0<=2; end
			5343: begin bcd3<=5;bcd2<=3;bcd1<=4;bcd0<=3; end
			5344: begin bcd3<=5;bcd2<=3;bcd1<=4;bcd0<=4; end
			5345: begin bcd3<=5;bcd2<=3;bcd1<=4;bcd0<=5; end
			5346: begin bcd3<=5;bcd2<=3;bcd1<=4;bcd0<=6; end
			5347: begin bcd3<=5;bcd2<=3;bcd1<=4;bcd0<=7; end
			5348: begin bcd3<=5;bcd2<=3;bcd1<=4;bcd0<=8; end
			5349: begin bcd3<=5;bcd2<=3;bcd1<=4;bcd0<=9; end
			5350: begin bcd3<=5;bcd2<=3;bcd1<=5;bcd0<=0; end
			5351: begin bcd3<=5;bcd2<=3;bcd1<=5;bcd0<=1; end
			5352: begin bcd3<=5;bcd2<=3;bcd1<=5;bcd0<=2; end
			5353: begin bcd3<=5;bcd2<=3;bcd1<=5;bcd0<=3; end
			5354: begin bcd3<=5;bcd2<=3;bcd1<=5;bcd0<=4; end
			5355: begin bcd3<=5;bcd2<=3;bcd1<=5;bcd0<=5; end
			5356: begin bcd3<=5;bcd2<=3;bcd1<=5;bcd0<=6; end
			5357: begin bcd3<=5;bcd2<=3;bcd1<=5;bcd0<=7; end
			5358: begin bcd3<=5;bcd2<=3;bcd1<=5;bcd0<=8; end
			5359: begin bcd3<=5;bcd2<=3;bcd1<=5;bcd0<=9; end
			5360: begin bcd3<=5;bcd2<=3;bcd1<=6;bcd0<=0; end
			5361: begin bcd3<=5;bcd2<=3;bcd1<=6;bcd0<=1; end
			5362: begin bcd3<=5;bcd2<=3;bcd1<=6;bcd0<=2; end
			5363: begin bcd3<=5;bcd2<=3;bcd1<=6;bcd0<=3; end
			5364: begin bcd3<=5;bcd2<=3;bcd1<=6;bcd0<=4; end
			5365: begin bcd3<=5;bcd2<=3;bcd1<=6;bcd0<=5; end
			5366: begin bcd3<=5;bcd2<=3;bcd1<=6;bcd0<=6; end
			5367: begin bcd3<=5;bcd2<=3;bcd1<=6;bcd0<=7; end
			5368: begin bcd3<=5;bcd2<=3;bcd1<=6;bcd0<=8; end
			5369: begin bcd3<=5;bcd2<=3;bcd1<=6;bcd0<=9; end
			5370: begin bcd3<=5;bcd2<=3;bcd1<=7;bcd0<=0; end
			5371: begin bcd3<=5;bcd2<=3;bcd1<=7;bcd0<=1; end
			5372: begin bcd3<=5;bcd2<=3;bcd1<=7;bcd0<=2; end
			5373: begin bcd3<=5;bcd2<=3;bcd1<=7;bcd0<=3; end
			5374: begin bcd3<=5;bcd2<=3;bcd1<=7;bcd0<=4; end
			5375: begin bcd3<=5;bcd2<=3;bcd1<=7;bcd0<=5; end
			5376: begin bcd3<=5;bcd2<=3;bcd1<=7;bcd0<=6; end
			5377: begin bcd3<=5;bcd2<=3;bcd1<=7;bcd0<=7; end
			5378: begin bcd3<=5;bcd2<=3;bcd1<=7;bcd0<=8; end
			5379: begin bcd3<=5;bcd2<=3;bcd1<=7;bcd0<=9; end
			5380: begin bcd3<=5;bcd2<=3;bcd1<=8;bcd0<=0; end
			5381: begin bcd3<=5;bcd2<=3;bcd1<=8;bcd0<=1; end
			5382: begin bcd3<=5;bcd2<=3;bcd1<=8;bcd0<=2; end
			5383: begin bcd3<=5;bcd2<=3;bcd1<=8;bcd0<=3; end
			5384: begin bcd3<=5;bcd2<=3;bcd1<=8;bcd0<=4; end
			5385: begin bcd3<=5;bcd2<=3;bcd1<=8;bcd0<=5; end
			5386: begin bcd3<=5;bcd2<=3;bcd1<=8;bcd0<=6; end
			5387: begin bcd3<=5;bcd2<=3;bcd1<=8;bcd0<=7; end
			5388: begin bcd3<=5;bcd2<=3;bcd1<=8;bcd0<=8; end
			5389: begin bcd3<=5;bcd2<=3;bcd1<=8;bcd0<=9; end
			5390: begin bcd3<=5;bcd2<=3;bcd1<=9;bcd0<=0; end
			5391: begin bcd3<=5;bcd2<=3;bcd1<=9;bcd0<=1; end
			5392: begin bcd3<=5;bcd2<=3;bcd1<=9;bcd0<=2; end
			5393: begin bcd3<=5;bcd2<=3;bcd1<=9;bcd0<=3; end
			5394: begin bcd3<=5;bcd2<=3;bcd1<=9;bcd0<=4; end
			5395: begin bcd3<=5;bcd2<=3;bcd1<=9;bcd0<=5; end
			5396: begin bcd3<=5;bcd2<=3;bcd1<=9;bcd0<=6; end
			5397: begin bcd3<=5;bcd2<=3;bcd1<=9;bcd0<=7; end
			5398: begin bcd3<=5;bcd2<=3;bcd1<=9;bcd0<=8; end
			5399: begin bcd3<=5;bcd2<=3;bcd1<=9;bcd0<=9; end
			5400: begin bcd3<=5;bcd2<=4;bcd1<=0;bcd0<=0; end
			5401: begin bcd3<=5;bcd2<=4;bcd1<=0;bcd0<=1; end
			5402: begin bcd3<=5;bcd2<=4;bcd1<=0;bcd0<=2; end
			5403: begin bcd3<=5;bcd2<=4;bcd1<=0;bcd0<=3; end
			5404: begin bcd3<=5;bcd2<=4;bcd1<=0;bcd0<=4; end
			5405: begin bcd3<=5;bcd2<=4;bcd1<=0;bcd0<=5; end
			5406: begin bcd3<=5;bcd2<=4;bcd1<=0;bcd0<=6; end
			5407: begin bcd3<=5;bcd2<=4;bcd1<=0;bcd0<=7; end
			5408: begin bcd3<=5;bcd2<=4;bcd1<=0;bcd0<=8; end
			5409: begin bcd3<=5;bcd2<=4;bcd1<=0;bcd0<=9; end
			5410: begin bcd3<=5;bcd2<=4;bcd1<=1;bcd0<=0; end
			5411: begin bcd3<=5;bcd2<=4;bcd1<=1;bcd0<=1; end
			5412: begin bcd3<=5;bcd2<=4;bcd1<=1;bcd0<=2; end
			5413: begin bcd3<=5;bcd2<=4;bcd1<=1;bcd0<=3; end
			5414: begin bcd3<=5;bcd2<=4;bcd1<=1;bcd0<=4; end
			5415: begin bcd3<=5;bcd2<=4;bcd1<=1;bcd0<=5; end
			5416: begin bcd3<=5;bcd2<=4;bcd1<=1;bcd0<=6; end
			5417: begin bcd3<=5;bcd2<=4;bcd1<=1;bcd0<=7; end
			5418: begin bcd3<=5;bcd2<=4;bcd1<=1;bcd0<=8; end
			5419: begin bcd3<=5;bcd2<=4;bcd1<=1;bcd0<=9; end
			5420: begin bcd3<=5;bcd2<=4;bcd1<=2;bcd0<=0; end
			5421: begin bcd3<=5;bcd2<=4;bcd1<=2;bcd0<=1; end
			5422: begin bcd3<=5;bcd2<=4;bcd1<=2;bcd0<=2; end
			5423: begin bcd3<=5;bcd2<=4;bcd1<=2;bcd0<=3; end
			5424: begin bcd3<=5;bcd2<=4;bcd1<=2;bcd0<=4; end
			5425: begin bcd3<=5;bcd2<=4;bcd1<=2;bcd0<=5; end
			5426: begin bcd3<=5;bcd2<=4;bcd1<=2;bcd0<=6; end
			5427: begin bcd3<=5;bcd2<=4;bcd1<=2;bcd0<=7; end
			5428: begin bcd3<=5;bcd2<=4;bcd1<=2;bcd0<=8; end
			5429: begin bcd3<=5;bcd2<=4;bcd1<=2;bcd0<=9; end
			5430: begin bcd3<=5;bcd2<=4;bcd1<=3;bcd0<=0; end
			5431: begin bcd3<=5;bcd2<=4;bcd1<=3;bcd0<=1; end
			5432: begin bcd3<=5;bcd2<=4;bcd1<=3;bcd0<=2; end
			5433: begin bcd3<=5;bcd2<=4;bcd1<=3;bcd0<=3; end
			5434: begin bcd3<=5;bcd2<=4;bcd1<=3;bcd0<=4; end
			5435: begin bcd3<=5;bcd2<=4;bcd1<=3;bcd0<=5; end
			5436: begin bcd3<=5;bcd2<=4;bcd1<=3;bcd0<=6; end
			5437: begin bcd3<=5;bcd2<=4;bcd1<=3;bcd0<=7; end
			5438: begin bcd3<=5;bcd2<=4;bcd1<=3;bcd0<=8; end
			5439: begin bcd3<=5;bcd2<=4;bcd1<=3;bcd0<=9; end
			5440: begin bcd3<=5;bcd2<=4;bcd1<=4;bcd0<=0; end
			5441: begin bcd3<=5;bcd2<=4;bcd1<=4;bcd0<=1; end
			5442: begin bcd3<=5;bcd2<=4;bcd1<=4;bcd0<=2; end
			5443: begin bcd3<=5;bcd2<=4;bcd1<=4;bcd0<=3; end
			5444: begin bcd3<=5;bcd2<=4;bcd1<=4;bcd0<=4; end
			5445: begin bcd3<=5;bcd2<=4;bcd1<=4;bcd0<=5; end
			5446: begin bcd3<=5;bcd2<=4;bcd1<=4;bcd0<=6; end
			5447: begin bcd3<=5;bcd2<=4;bcd1<=4;bcd0<=7; end
			5448: begin bcd3<=5;bcd2<=4;bcd1<=4;bcd0<=8; end
			5449: begin bcd3<=5;bcd2<=4;bcd1<=4;bcd0<=9; end
			5450: begin bcd3<=5;bcd2<=4;bcd1<=5;bcd0<=0; end
			5451: begin bcd3<=5;bcd2<=4;bcd1<=5;bcd0<=1; end
			5452: begin bcd3<=5;bcd2<=4;bcd1<=5;bcd0<=2; end
			5453: begin bcd3<=5;bcd2<=4;bcd1<=5;bcd0<=3; end
			5454: begin bcd3<=5;bcd2<=4;bcd1<=5;bcd0<=4; end
			5455: begin bcd3<=5;bcd2<=4;bcd1<=5;bcd0<=5; end
			5456: begin bcd3<=5;bcd2<=4;bcd1<=5;bcd0<=6; end
			5457: begin bcd3<=5;bcd2<=4;bcd1<=5;bcd0<=7; end
			5458: begin bcd3<=5;bcd2<=4;bcd1<=5;bcd0<=8; end
			5459: begin bcd3<=5;bcd2<=4;bcd1<=5;bcd0<=9; end
			5460: begin bcd3<=5;bcd2<=4;bcd1<=6;bcd0<=0; end
			5461: begin bcd3<=5;bcd2<=4;bcd1<=6;bcd0<=1; end
			5462: begin bcd3<=5;bcd2<=4;bcd1<=6;bcd0<=2; end
			5463: begin bcd3<=5;bcd2<=4;bcd1<=6;bcd0<=3; end
			5464: begin bcd3<=5;bcd2<=4;bcd1<=6;bcd0<=4; end
			5465: begin bcd3<=5;bcd2<=4;bcd1<=6;bcd0<=5; end
			5466: begin bcd3<=5;bcd2<=4;bcd1<=6;bcd0<=6; end
			5467: begin bcd3<=5;bcd2<=4;bcd1<=6;bcd0<=7; end
			5468: begin bcd3<=5;bcd2<=4;bcd1<=6;bcd0<=8; end
			5469: begin bcd3<=5;bcd2<=4;bcd1<=6;bcd0<=9; end
			5470: begin bcd3<=5;bcd2<=4;bcd1<=7;bcd0<=0; end
			5471: begin bcd3<=5;bcd2<=4;bcd1<=7;bcd0<=1; end
			5472: begin bcd3<=5;bcd2<=4;bcd1<=7;bcd0<=2; end
			5473: begin bcd3<=5;bcd2<=4;bcd1<=7;bcd0<=3; end
			5474: begin bcd3<=5;bcd2<=4;bcd1<=7;bcd0<=4; end
			5475: begin bcd3<=5;bcd2<=4;bcd1<=7;bcd0<=5; end
			5476: begin bcd3<=5;bcd2<=4;bcd1<=7;bcd0<=6; end
			5477: begin bcd3<=5;bcd2<=4;bcd1<=7;bcd0<=7; end
			5478: begin bcd3<=5;bcd2<=4;bcd1<=7;bcd0<=8; end
			5479: begin bcd3<=5;bcd2<=4;bcd1<=7;bcd0<=9; end
			5480: begin bcd3<=5;bcd2<=4;bcd1<=8;bcd0<=0; end
			5481: begin bcd3<=5;bcd2<=4;bcd1<=8;bcd0<=1; end
			5482: begin bcd3<=5;bcd2<=4;bcd1<=8;bcd0<=2; end
			5483: begin bcd3<=5;bcd2<=4;bcd1<=8;bcd0<=3; end
			5484: begin bcd3<=5;bcd2<=4;bcd1<=8;bcd0<=4; end
			5485: begin bcd3<=5;bcd2<=4;bcd1<=8;bcd0<=5; end
			5486: begin bcd3<=5;bcd2<=4;bcd1<=8;bcd0<=6; end
			5487: begin bcd3<=5;bcd2<=4;bcd1<=8;bcd0<=7; end
			5488: begin bcd3<=5;bcd2<=4;bcd1<=8;bcd0<=8; end
			5489: begin bcd3<=5;bcd2<=4;bcd1<=8;bcd0<=9; end
			5490: begin bcd3<=5;bcd2<=4;bcd1<=9;bcd0<=0; end
			5491: begin bcd3<=5;bcd2<=4;bcd1<=9;bcd0<=1; end
			5492: begin bcd3<=5;bcd2<=4;bcd1<=9;bcd0<=2; end
			5493: begin bcd3<=5;bcd2<=4;bcd1<=9;bcd0<=3; end
			5494: begin bcd3<=5;bcd2<=4;bcd1<=9;bcd0<=4; end
			5495: begin bcd3<=5;bcd2<=4;bcd1<=9;bcd0<=5; end
			5496: begin bcd3<=5;bcd2<=4;bcd1<=9;bcd0<=6; end
			5497: begin bcd3<=5;bcd2<=4;bcd1<=9;bcd0<=7; end
			5498: begin bcd3<=5;bcd2<=4;bcd1<=9;bcd0<=8; end
			5499: begin bcd3<=5;bcd2<=4;bcd1<=9;bcd0<=9; end
			5500: begin bcd3<=5;bcd2<=5;bcd1<=0;bcd0<=0; end
			5501: begin bcd3<=5;bcd2<=5;bcd1<=0;bcd0<=1; end
			5502: begin bcd3<=5;bcd2<=5;bcd1<=0;bcd0<=2; end
			5503: begin bcd3<=5;bcd2<=5;bcd1<=0;bcd0<=3; end
			5504: begin bcd3<=5;bcd2<=5;bcd1<=0;bcd0<=4; end
			5505: begin bcd3<=5;bcd2<=5;bcd1<=0;bcd0<=5; end
			5506: begin bcd3<=5;bcd2<=5;bcd1<=0;bcd0<=6; end
			5507: begin bcd3<=5;bcd2<=5;bcd1<=0;bcd0<=7; end
			5508: begin bcd3<=5;bcd2<=5;bcd1<=0;bcd0<=8; end
			5509: begin bcd3<=5;bcd2<=5;bcd1<=0;bcd0<=9; end
			5510: begin bcd3<=5;bcd2<=5;bcd1<=1;bcd0<=0; end
			5511: begin bcd3<=5;bcd2<=5;bcd1<=1;bcd0<=1; end
			5512: begin bcd3<=5;bcd2<=5;bcd1<=1;bcd0<=2; end
			5513: begin bcd3<=5;bcd2<=5;bcd1<=1;bcd0<=3; end
			5514: begin bcd3<=5;bcd2<=5;bcd1<=1;bcd0<=4; end
			5515: begin bcd3<=5;bcd2<=5;bcd1<=1;bcd0<=5; end
			5516: begin bcd3<=5;bcd2<=5;bcd1<=1;bcd0<=6; end
			5517: begin bcd3<=5;bcd2<=5;bcd1<=1;bcd0<=7; end
			5518: begin bcd3<=5;bcd2<=5;bcd1<=1;bcd0<=8; end
			5519: begin bcd3<=5;bcd2<=5;bcd1<=1;bcd0<=9; end
			5520: begin bcd3<=5;bcd2<=5;bcd1<=2;bcd0<=0; end
			5521: begin bcd3<=5;bcd2<=5;bcd1<=2;bcd0<=1; end
			5522: begin bcd3<=5;bcd2<=5;bcd1<=2;bcd0<=2; end
			5523: begin bcd3<=5;bcd2<=5;bcd1<=2;bcd0<=3; end
			5524: begin bcd3<=5;bcd2<=5;bcd1<=2;bcd0<=4; end
			5525: begin bcd3<=5;bcd2<=5;bcd1<=2;bcd0<=5; end
			5526: begin bcd3<=5;bcd2<=5;bcd1<=2;bcd0<=6; end
			5527: begin bcd3<=5;bcd2<=5;bcd1<=2;bcd0<=7; end
			5528: begin bcd3<=5;bcd2<=5;bcd1<=2;bcd0<=8; end
			5529: begin bcd3<=5;bcd2<=5;bcd1<=2;bcd0<=9; end
			5530: begin bcd3<=5;bcd2<=5;bcd1<=3;bcd0<=0; end
			5531: begin bcd3<=5;bcd2<=5;bcd1<=3;bcd0<=1; end
			5532: begin bcd3<=5;bcd2<=5;bcd1<=3;bcd0<=2; end
			5533: begin bcd3<=5;bcd2<=5;bcd1<=3;bcd0<=3; end
			5534: begin bcd3<=5;bcd2<=5;bcd1<=3;bcd0<=4; end
			5535: begin bcd3<=5;bcd2<=5;bcd1<=3;bcd0<=5; end
			5536: begin bcd3<=5;bcd2<=5;bcd1<=3;bcd0<=6; end
			5537: begin bcd3<=5;bcd2<=5;bcd1<=3;bcd0<=7; end
			5538: begin bcd3<=5;bcd2<=5;bcd1<=3;bcd0<=8; end
			5539: begin bcd3<=5;bcd2<=5;bcd1<=3;bcd0<=9; end
			5540: begin bcd3<=5;bcd2<=5;bcd1<=4;bcd0<=0; end
			5541: begin bcd3<=5;bcd2<=5;bcd1<=4;bcd0<=1; end
			5542: begin bcd3<=5;bcd2<=5;bcd1<=4;bcd0<=2; end
			5543: begin bcd3<=5;bcd2<=5;bcd1<=4;bcd0<=3; end
			5544: begin bcd3<=5;bcd2<=5;bcd1<=4;bcd0<=4; end
			5545: begin bcd3<=5;bcd2<=5;bcd1<=4;bcd0<=5; end
			5546: begin bcd3<=5;bcd2<=5;bcd1<=4;bcd0<=6; end
			5547: begin bcd3<=5;bcd2<=5;bcd1<=4;bcd0<=7; end
			5548: begin bcd3<=5;bcd2<=5;bcd1<=4;bcd0<=8; end
			5549: begin bcd3<=5;bcd2<=5;bcd1<=4;bcd0<=9; end
			5550: begin bcd3<=5;bcd2<=5;bcd1<=5;bcd0<=0; end
			5551: begin bcd3<=5;bcd2<=5;bcd1<=5;bcd0<=1; end
			5552: begin bcd3<=5;bcd2<=5;bcd1<=5;bcd0<=2; end
			5553: begin bcd3<=5;bcd2<=5;bcd1<=5;bcd0<=3; end
			5554: begin bcd3<=5;bcd2<=5;bcd1<=5;bcd0<=4; end
			5555: begin bcd3<=5;bcd2<=5;bcd1<=5;bcd0<=5; end
			5556: begin bcd3<=5;bcd2<=5;bcd1<=5;bcd0<=6; end
			5557: begin bcd3<=5;bcd2<=5;bcd1<=5;bcd0<=7; end
			5558: begin bcd3<=5;bcd2<=5;bcd1<=5;bcd0<=8; end
			5559: begin bcd3<=5;bcd2<=5;bcd1<=5;bcd0<=9; end
			5560: begin bcd3<=5;bcd2<=5;bcd1<=6;bcd0<=0; end
			5561: begin bcd3<=5;bcd2<=5;bcd1<=6;bcd0<=1; end
			5562: begin bcd3<=5;bcd2<=5;bcd1<=6;bcd0<=2; end
			5563: begin bcd3<=5;bcd2<=5;bcd1<=6;bcd0<=3; end
			5564: begin bcd3<=5;bcd2<=5;bcd1<=6;bcd0<=4; end
			5565: begin bcd3<=5;bcd2<=5;bcd1<=6;bcd0<=5; end
			5566: begin bcd3<=5;bcd2<=5;bcd1<=6;bcd0<=6; end
			5567: begin bcd3<=5;bcd2<=5;bcd1<=6;bcd0<=7; end
			5568: begin bcd3<=5;bcd2<=5;bcd1<=6;bcd0<=8; end
			5569: begin bcd3<=5;bcd2<=5;bcd1<=6;bcd0<=9; end
			5570: begin bcd3<=5;bcd2<=5;bcd1<=7;bcd0<=0; end
			5571: begin bcd3<=5;bcd2<=5;bcd1<=7;bcd0<=1; end
			5572: begin bcd3<=5;bcd2<=5;bcd1<=7;bcd0<=2; end
			5573: begin bcd3<=5;bcd2<=5;bcd1<=7;bcd0<=3; end
			5574: begin bcd3<=5;bcd2<=5;bcd1<=7;bcd0<=4; end
			5575: begin bcd3<=5;bcd2<=5;bcd1<=7;bcd0<=5; end
			5576: begin bcd3<=5;bcd2<=5;bcd1<=7;bcd0<=6; end
			5577: begin bcd3<=5;bcd2<=5;bcd1<=7;bcd0<=7; end
			5578: begin bcd3<=5;bcd2<=5;bcd1<=7;bcd0<=8; end
			5579: begin bcd3<=5;bcd2<=5;bcd1<=7;bcd0<=9; end
			5580: begin bcd3<=5;bcd2<=5;bcd1<=8;bcd0<=0; end
			5581: begin bcd3<=5;bcd2<=5;bcd1<=8;bcd0<=1; end
			5582: begin bcd3<=5;bcd2<=5;bcd1<=8;bcd0<=2; end
			5583: begin bcd3<=5;bcd2<=5;bcd1<=8;bcd0<=3; end
			5584: begin bcd3<=5;bcd2<=5;bcd1<=8;bcd0<=4; end
			5585: begin bcd3<=5;bcd2<=5;bcd1<=8;bcd0<=5; end
			5586: begin bcd3<=5;bcd2<=5;bcd1<=8;bcd0<=6; end
			5587: begin bcd3<=5;bcd2<=5;bcd1<=8;bcd0<=7; end
			5588: begin bcd3<=5;bcd2<=5;bcd1<=8;bcd0<=8; end
			5589: begin bcd3<=5;bcd2<=5;bcd1<=8;bcd0<=9; end
			5590: begin bcd3<=5;bcd2<=5;bcd1<=9;bcd0<=0; end
			5591: begin bcd3<=5;bcd2<=5;bcd1<=9;bcd0<=1; end
			5592: begin bcd3<=5;bcd2<=5;bcd1<=9;bcd0<=2; end
			5593: begin bcd3<=5;bcd2<=5;bcd1<=9;bcd0<=3; end
			5594: begin bcd3<=5;bcd2<=5;bcd1<=9;bcd0<=4; end
			5595: begin bcd3<=5;bcd2<=5;bcd1<=9;bcd0<=5; end
			5596: begin bcd3<=5;bcd2<=5;bcd1<=9;bcd0<=6; end
			5597: begin bcd3<=5;bcd2<=5;bcd1<=9;bcd0<=7; end
			5598: begin bcd3<=5;bcd2<=5;bcd1<=9;bcd0<=8; end
			5599: begin bcd3<=5;bcd2<=5;bcd1<=9;bcd0<=9; end
			5600: begin bcd3<=5;bcd2<=6;bcd1<=0;bcd0<=0; end
			5601: begin bcd3<=5;bcd2<=6;bcd1<=0;bcd0<=1; end
			5602: begin bcd3<=5;bcd2<=6;bcd1<=0;bcd0<=2; end
			5603: begin bcd3<=5;bcd2<=6;bcd1<=0;bcd0<=3; end
			5604: begin bcd3<=5;bcd2<=6;bcd1<=0;bcd0<=4; end
			5605: begin bcd3<=5;bcd2<=6;bcd1<=0;bcd0<=5; end
			5606: begin bcd3<=5;bcd2<=6;bcd1<=0;bcd0<=6; end
			5607: begin bcd3<=5;bcd2<=6;bcd1<=0;bcd0<=7; end
			5608: begin bcd3<=5;bcd2<=6;bcd1<=0;bcd0<=8; end
			5609: begin bcd3<=5;bcd2<=6;bcd1<=0;bcd0<=9; end
			5610: begin bcd3<=5;bcd2<=6;bcd1<=1;bcd0<=0; end
			5611: begin bcd3<=5;bcd2<=6;bcd1<=1;bcd0<=1; end
			5612: begin bcd3<=5;bcd2<=6;bcd1<=1;bcd0<=2; end
			5613: begin bcd3<=5;bcd2<=6;bcd1<=1;bcd0<=3; end
			5614: begin bcd3<=5;bcd2<=6;bcd1<=1;bcd0<=4; end
			5615: begin bcd3<=5;bcd2<=6;bcd1<=1;bcd0<=5; end
			5616: begin bcd3<=5;bcd2<=6;bcd1<=1;bcd0<=6; end
			5617: begin bcd3<=5;bcd2<=6;bcd1<=1;bcd0<=7; end
			5618: begin bcd3<=5;bcd2<=6;bcd1<=1;bcd0<=8; end
			5619: begin bcd3<=5;bcd2<=6;bcd1<=1;bcd0<=9; end
			5620: begin bcd3<=5;bcd2<=6;bcd1<=2;bcd0<=0; end
			5621: begin bcd3<=5;bcd2<=6;bcd1<=2;bcd0<=1; end
			5622: begin bcd3<=5;bcd2<=6;bcd1<=2;bcd0<=2; end
			5623: begin bcd3<=5;bcd2<=6;bcd1<=2;bcd0<=3; end
			5624: begin bcd3<=5;bcd2<=6;bcd1<=2;bcd0<=4; end
			5625: begin bcd3<=5;bcd2<=6;bcd1<=2;bcd0<=5; end
			5626: begin bcd3<=5;bcd2<=6;bcd1<=2;bcd0<=6; end
			5627: begin bcd3<=5;bcd2<=6;bcd1<=2;bcd0<=7; end
			5628: begin bcd3<=5;bcd2<=6;bcd1<=2;bcd0<=8; end
			5629: begin bcd3<=5;bcd2<=6;bcd1<=2;bcd0<=9; end
			5630: begin bcd3<=5;bcd2<=6;bcd1<=3;bcd0<=0; end
			5631: begin bcd3<=5;bcd2<=6;bcd1<=3;bcd0<=1; end
			5632: begin bcd3<=5;bcd2<=6;bcd1<=3;bcd0<=2; end
			5633: begin bcd3<=5;bcd2<=6;bcd1<=3;bcd0<=3; end
			5634: begin bcd3<=5;bcd2<=6;bcd1<=3;bcd0<=4; end
			5635: begin bcd3<=5;bcd2<=6;bcd1<=3;bcd0<=5; end
			5636: begin bcd3<=5;bcd2<=6;bcd1<=3;bcd0<=6; end
			5637: begin bcd3<=5;bcd2<=6;bcd1<=3;bcd0<=7; end
			5638: begin bcd3<=5;bcd2<=6;bcd1<=3;bcd0<=8; end
			5639: begin bcd3<=5;bcd2<=6;bcd1<=3;bcd0<=9; end
			5640: begin bcd3<=5;bcd2<=6;bcd1<=4;bcd0<=0; end
			5641: begin bcd3<=5;bcd2<=6;bcd1<=4;bcd0<=1; end
			5642: begin bcd3<=5;bcd2<=6;bcd1<=4;bcd0<=2; end
			5643: begin bcd3<=5;bcd2<=6;bcd1<=4;bcd0<=3; end
			5644: begin bcd3<=5;bcd2<=6;bcd1<=4;bcd0<=4; end
			5645: begin bcd3<=5;bcd2<=6;bcd1<=4;bcd0<=5; end
			5646: begin bcd3<=5;bcd2<=6;bcd1<=4;bcd0<=6; end
			5647: begin bcd3<=5;bcd2<=6;bcd1<=4;bcd0<=7; end
			5648: begin bcd3<=5;bcd2<=6;bcd1<=4;bcd0<=8; end
			5649: begin bcd3<=5;bcd2<=6;bcd1<=4;bcd0<=9; end
			5650: begin bcd3<=5;bcd2<=6;bcd1<=5;bcd0<=0; end
			5651: begin bcd3<=5;bcd2<=6;bcd1<=5;bcd0<=1; end
			5652: begin bcd3<=5;bcd2<=6;bcd1<=5;bcd0<=2; end
			5653: begin bcd3<=5;bcd2<=6;bcd1<=5;bcd0<=3; end
			5654: begin bcd3<=5;bcd2<=6;bcd1<=5;bcd0<=4; end
			5655: begin bcd3<=5;bcd2<=6;bcd1<=5;bcd0<=5; end
			5656: begin bcd3<=5;bcd2<=6;bcd1<=5;bcd0<=6; end
			5657: begin bcd3<=5;bcd2<=6;bcd1<=5;bcd0<=7; end
			5658: begin bcd3<=5;bcd2<=6;bcd1<=5;bcd0<=8; end
			5659: begin bcd3<=5;bcd2<=6;bcd1<=5;bcd0<=9; end
			5660: begin bcd3<=5;bcd2<=6;bcd1<=6;bcd0<=0; end
			5661: begin bcd3<=5;bcd2<=6;bcd1<=6;bcd0<=1; end
			5662: begin bcd3<=5;bcd2<=6;bcd1<=6;bcd0<=2; end
			5663: begin bcd3<=5;bcd2<=6;bcd1<=6;bcd0<=3; end
			5664: begin bcd3<=5;bcd2<=6;bcd1<=6;bcd0<=4; end
			5665: begin bcd3<=5;bcd2<=6;bcd1<=6;bcd0<=5; end
			5666: begin bcd3<=5;bcd2<=6;bcd1<=6;bcd0<=6; end
			5667: begin bcd3<=5;bcd2<=6;bcd1<=6;bcd0<=7; end
			5668: begin bcd3<=5;bcd2<=6;bcd1<=6;bcd0<=8; end
			5669: begin bcd3<=5;bcd2<=6;bcd1<=6;bcd0<=9; end
			5670: begin bcd3<=5;bcd2<=6;bcd1<=7;bcd0<=0; end
			5671: begin bcd3<=5;bcd2<=6;bcd1<=7;bcd0<=1; end
			5672: begin bcd3<=5;bcd2<=6;bcd1<=7;bcd0<=2; end
			5673: begin bcd3<=5;bcd2<=6;bcd1<=7;bcd0<=3; end
			5674: begin bcd3<=5;bcd2<=6;bcd1<=7;bcd0<=4; end
			5675: begin bcd3<=5;bcd2<=6;bcd1<=7;bcd0<=5; end
			5676: begin bcd3<=5;bcd2<=6;bcd1<=7;bcd0<=6; end
			5677: begin bcd3<=5;bcd2<=6;bcd1<=7;bcd0<=7; end
			5678: begin bcd3<=5;bcd2<=6;bcd1<=7;bcd0<=8; end
			5679: begin bcd3<=5;bcd2<=6;bcd1<=7;bcd0<=9; end
			5680: begin bcd3<=5;bcd2<=6;bcd1<=8;bcd0<=0; end
			5681: begin bcd3<=5;bcd2<=6;bcd1<=8;bcd0<=1; end
			5682: begin bcd3<=5;bcd2<=6;bcd1<=8;bcd0<=2; end
			5683: begin bcd3<=5;bcd2<=6;bcd1<=8;bcd0<=3; end
			5684: begin bcd3<=5;bcd2<=6;bcd1<=8;bcd0<=4; end
			5685: begin bcd3<=5;bcd2<=6;bcd1<=8;bcd0<=5; end
			5686: begin bcd3<=5;bcd2<=6;bcd1<=8;bcd0<=6; end
			5687: begin bcd3<=5;bcd2<=6;bcd1<=8;bcd0<=7; end
			5688: begin bcd3<=5;bcd2<=6;bcd1<=8;bcd0<=8; end
			5689: begin bcd3<=5;bcd2<=6;bcd1<=8;bcd0<=9; end
			5690: begin bcd3<=5;bcd2<=6;bcd1<=9;bcd0<=0; end
			5691: begin bcd3<=5;bcd2<=6;bcd1<=9;bcd0<=1; end
			5692: begin bcd3<=5;bcd2<=6;bcd1<=9;bcd0<=2; end
			5693: begin bcd3<=5;bcd2<=6;bcd1<=9;bcd0<=3; end
			5694: begin bcd3<=5;bcd2<=6;bcd1<=9;bcd0<=4; end
			5695: begin bcd3<=5;bcd2<=6;bcd1<=9;bcd0<=5; end
			5696: begin bcd3<=5;bcd2<=6;bcd1<=9;bcd0<=6; end
			5697: begin bcd3<=5;bcd2<=6;bcd1<=9;bcd0<=7; end
			5698: begin bcd3<=5;bcd2<=6;bcd1<=9;bcd0<=8; end
			5699: begin bcd3<=5;bcd2<=6;bcd1<=9;bcd0<=9; end
			5700: begin bcd3<=5;bcd2<=7;bcd1<=0;bcd0<=0; end
			5701: begin bcd3<=5;bcd2<=7;bcd1<=0;bcd0<=1; end
			5702: begin bcd3<=5;bcd2<=7;bcd1<=0;bcd0<=2; end
			5703: begin bcd3<=5;bcd2<=7;bcd1<=0;bcd0<=3; end
			5704: begin bcd3<=5;bcd2<=7;bcd1<=0;bcd0<=4; end
			5705: begin bcd3<=5;bcd2<=7;bcd1<=0;bcd0<=5; end
			5706: begin bcd3<=5;bcd2<=7;bcd1<=0;bcd0<=6; end
			5707: begin bcd3<=5;bcd2<=7;bcd1<=0;bcd0<=7; end
			5708: begin bcd3<=5;bcd2<=7;bcd1<=0;bcd0<=8; end
			5709: begin bcd3<=5;bcd2<=7;bcd1<=0;bcd0<=9; end
			5710: begin bcd3<=5;bcd2<=7;bcd1<=1;bcd0<=0; end
			5711: begin bcd3<=5;bcd2<=7;bcd1<=1;bcd0<=1; end
			5712: begin bcd3<=5;bcd2<=7;bcd1<=1;bcd0<=2; end
			5713: begin bcd3<=5;bcd2<=7;bcd1<=1;bcd0<=3; end
			5714: begin bcd3<=5;bcd2<=7;bcd1<=1;bcd0<=4; end
			5715: begin bcd3<=5;bcd2<=7;bcd1<=1;bcd0<=5; end
			5716: begin bcd3<=5;bcd2<=7;bcd1<=1;bcd0<=6; end
			5717: begin bcd3<=5;bcd2<=7;bcd1<=1;bcd0<=7; end
			5718: begin bcd3<=5;bcd2<=7;bcd1<=1;bcd0<=8; end
			5719: begin bcd3<=5;bcd2<=7;bcd1<=1;bcd0<=9; end
			5720: begin bcd3<=5;bcd2<=7;bcd1<=2;bcd0<=0; end
			5721: begin bcd3<=5;bcd2<=7;bcd1<=2;bcd0<=1; end
			5722: begin bcd3<=5;bcd2<=7;bcd1<=2;bcd0<=2; end
			5723: begin bcd3<=5;bcd2<=7;bcd1<=2;bcd0<=3; end
			5724: begin bcd3<=5;bcd2<=7;bcd1<=2;bcd0<=4; end
			5725: begin bcd3<=5;bcd2<=7;bcd1<=2;bcd0<=5; end
			5726: begin bcd3<=5;bcd2<=7;bcd1<=2;bcd0<=6; end
			5727: begin bcd3<=5;bcd2<=7;bcd1<=2;bcd0<=7; end
			5728: begin bcd3<=5;bcd2<=7;bcd1<=2;bcd0<=8; end
			5729: begin bcd3<=5;bcd2<=7;bcd1<=2;bcd0<=9; end
			5730: begin bcd3<=5;bcd2<=7;bcd1<=3;bcd0<=0; end
			5731: begin bcd3<=5;bcd2<=7;bcd1<=3;bcd0<=1; end
			5732: begin bcd3<=5;bcd2<=7;bcd1<=3;bcd0<=2; end
			5733: begin bcd3<=5;bcd2<=7;bcd1<=3;bcd0<=3; end
			5734: begin bcd3<=5;bcd2<=7;bcd1<=3;bcd0<=4; end
			5735: begin bcd3<=5;bcd2<=7;bcd1<=3;bcd0<=5; end
			5736: begin bcd3<=5;bcd2<=7;bcd1<=3;bcd0<=6; end
			5737: begin bcd3<=5;bcd2<=7;bcd1<=3;bcd0<=7; end
			5738: begin bcd3<=5;bcd2<=7;bcd1<=3;bcd0<=8; end
			5739: begin bcd3<=5;bcd2<=7;bcd1<=3;bcd0<=9; end
			5740: begin bcd3<=5;bcd2<=7;bcd1<=4;bcd0<=0; end
			5741: begin bcd3<=5;bcd2<=7;bcd1<=4;bcd0<=1; end
			5742: begin bcd3<=5;bcd2<=7;bcd1<=4;bcd0<=2; end
			5743: begin bcd3<=5;bcd2<=7;bcd1<=4;bcd0<=3; end
			5744: begin bcd3<=5;bcd2<=7;bcd1<=4;bcd0<=4; end
			5745: begin bcd3<=5;bcd2<=7;bcd1<=4;bcd0<=5; end
			5746: begin bcd3<=5;bcd2<=7;bcd1<=4;bcd0<=6; end
			5747: begin bcd3<=5;bcd2<=7;bcd1<=4;bcd0<=7; end
			5748: begin bcd3<=5;bcd2<=7;bcd1<=4;bcd0<=8; end
			5749: begin bcd3<=5;bcd2<=7;bcd1<=4;bcd0<=9; end
			5750: begin bcd3<=5;bcd2<=7;bcd1<=5;bcd0<=0; end
			5751: begin bcd3<=5;bcd2<=7;bcd1<=5;bcd0<=1; end
			5752: begin bcd3<=5;bcd2<=7;bcd1<=5;bcd0<=2; end
			5753: begin bcd3<=5;bcd2<=7;bcd1<=5;bcd0<=3; end
			5754: begin bcd3<=5;bcd2<=7;bcd1<=5;bcd0<=4; end
			5755: begin bcd3<=5;bcd2<=7;bcd1<=5;bcd0<=5; end
			5756: begin bcd3<=5;bcd2<=7;bcd1<=5;bcd0<=6; end
			5757: begin bcd3<=5;bcd2<=7;bcd1<=5;bcd0<=7; end
			5758: begin bcd3<=5;bcd2<=7;bcd1<=5;bcd0<=8; end
			5759: begin bcd3<=5;bcd2<=7;bcd1<=5;bcd0<=9; end
			5760: begin bcd3<=5;bcd2<=7;bcd1<=6;bcd0<=0; end
			5761: begin bcd3<=5;bcd2<=7;bcd1<=6;bcd0<=1; end
			5762: begin bcd3<=5;bcd2<=7;bcd1<=6;bcd0<=2; end
			5763: begin bcd3<=5;bcd2<=7;bcd1<=6;bcd0<=3; end
			5764: begin bcd3<=5;bcd2<=7;bcd1<=6;bcd0<=4; end
			5765: begin bcd3<=5;bcd2<=7;bcd1<=6;bcd0<=5; end
			5766: begin bcd3<=5;bcd2<=7;bcd1<=6;bcd0<=6; end
			5767: begin bcd3<=5;bcd2<=7;bcd1<=6;bcd0<=7; end
			5768: begin bcd3<=5;bcd2<=7;bcd1<=6;bcd0<=8; end
			5769: begin bcd3<=5;bcd2<=7;bcd1<=6;bcd0<=9; end
			5770: begin bcd3<=5;bcd2<=7;bcd1<=7;bcd0<=0; end
			5771: begin bcd3<=5;bcd2<=7;bcd1<=7;bcd0<=1; end
			5772: begin bcd3<=5;bcd2<=7;bcd1<=7;bcd0<=2; end
			5773: begin bcd3<=5;bcd2<=7;bcd1<=7;bcd0<=3; end
			5774: begin bcd3<=5;bcd2<=7;bcd1<=7;bcd0<=4; end
			5775: begin bcd3<=5;bcd2<=7;bcd1<=7;bcd0<=5; end
			5776: begin bcd3<=5;bcd2<=7;bcd1<=7;bcd0<=6; end
			5777: begin bcd3<=5;bcd2<=7;bcd1<=7;bcd0<=7; end
			5778: begin bcd3<=5;bcd2<=7;bcd1<=7;bcd0<=8; end
			5779: begin bcd3<=5;bcd2<=7;bcd1<=7;bcd0<=9; end
			5780: begin bcd3<=5;bcd2<=7;bcd1<=8;bcd0<=0; end
			5781: begin bcd3<=5;bcd2<=7;bcd1<=8;bcd0<=1; end
			5782: begin bcd3<=5;bcd2<=7;bcd1<=8;bcd0<=2; end
			5783: begin bcd3<=5;bcd2<=7;bcd1<=8;bcd0<=3; end
			5784: begin bcd3<=5;bcd2<=7;bcd1<=8;bcd0<=4; end
			5785: begin bcd3<=5;bcd2<=7;bcd1<=8;bcd0<=5; end
			5786: begin bcd3<=5;bcd2<=7;bcd1<=8;bcd0<=6; end
			5787: begin bcd3<=5;bcd2<=7;bcd1<=8;bcd0<=7; end
			5788: begin bcd3<=5;bcd2<=7;bcd1<=8;bcd0<=8; end
			5789: begin bcd3<=5;bcd2<=7;bcd1<=8;bcd0<=9; end
			5790: begin bcd3<=5;bcd2<=7;bcd1<=9;bcd0<=0; end
			5791: begin bcd3<=5;bcd2<=7;bcd1<=9;bcd0<=1; end
			5792: begin bcd3<=5;bcd2<=7;bcd1<=9;bcd0<=2; end
			5793: begin bcd3<=5;bcd2<=7;bcd1<=9;bcd0<=3; end
			5794: begin bcd3<=5;bcd2<=7;bcd1<=9;bcd0<=4; end
			5795: begin bcd3<=5;bcd2<=7;bcd1<=9;bcd0<=5; end
			5796: begin bcd3<=5;bcd2<=7;bcd1<=9;bcd0<=6; end
			5797: begin bcd3<=5;bcd2<=7;bcd1<=9;bcd0<=7; end
			5798: begin bcd3<=5;bcd2<=7;bcd1<=9;bcd0<=8; end
			5799: begin bcd3<=5;bcd2<=7;bcd1<=9;bcd0<=9; end
			5800: begin bcd3<=5;bcd2<=8;bcd1<=0;bcd0<=0; end
			5801: begin bcd3<=5;bcd2<=8;bcd1<=0;bcd0<=1; end
			5802: begin bcd3<=5;bcd2<=8;bcd1<=0;bcd0<=2; end
			5803: begin bcd3<=5;bcd2<=8;bcd1<=0;bcd0<=3; end
			5804: begin bcd3<=5;bcd2<=8;bcd1<=0;bcd0<=4; end
			5805: begin bcd3<=5;bcd2<=8;bcd1<=0;bcd0<=5; end
			5806: begin bcd3<=5;bcd2<=8;bcd1<=0;bcd0<=6; end
			5807: begin bcd3<=5;bcd2<=8;bcd1<=0;bcd0<=7; end
			5808: begin bcd3<=5;bcd2<=8;bcd1<=0;bcd0<=8; end
			5809: begin bcd3<=5;bcd2<=8;bcd1<=0;bcd0<=9; end
			5810: begin bcd3<=5;bcd2<=8;bcd1<=1;bcd0<=0; end
			5811: begin bcd3<=5;bcd2<=8;bcd1<=1;bcd0<=1; end
			5812: begin bcd3<=5;bcd2<=8;bcd1<=1;bcd0<=2; end
			5813: begin bcd3<=5;bcd2<=8;bcd1<=1;bcd0<=3; end
			5814: begin bcd3<=5;bcd2<=8;bcd1<=1;bcd0<=4; end
			5815: begin bcd3<=5;bcd2<=8;bcd1<=1;bcd0<=5; end
			5816: begin bcd3<=5;bcd2<=8;bcd1<=1;bcd0<=6; end
			5817: begin bcd3<=5;bcd2<=8;bcd1<=1;bcd0<=7; end
			5818: begin bcd3<=5;bcd2<=8;bcd1<=1;bcd0<=8; end
			5819: begin bcd3<=5;bcd2<=8;bcd1<=1;bcd0<=9; end
			5820: begin bcd3<=5;bcd2<=8;bcd1<=2;bcd0<=0; end
			5821: begin bcd3<=5;bcd2<=8;bcd1<=2;bcd0<=1; end
			5822: begin bcd3<=5;bcd2<=8;bcd1<=2;bcd0<=2; end
			5823: begin bcd3<=5;bcd2<=8;bcd1<=2;bcd0<=3; end
			5824: begin bcd3<=5;bcd2<=8;bcd1<=2;bcd0<=4; end
			5825: begin bcd3<=5;bcd2<=8;bcd1<=2;bcd0<=5; end
			5826: begin bcd3<=5;bcd2<=8;bcd1<=2;bcd0<=6; end
			5827: begin bcd3<=5;bcd2<=8;bcd1<=2;bcd0<=7; end
			5828: begin bcd3<=5;bcd2<=8;bcd1<=2;bcd0<=8; end
			5829: begin bcd3<=5;bcd2<=8;bcd1<=2;bcd0<=9; end
			5830: begin bcd3<=5;bcd2<=8;bcd1<=3;bcd0<=0; end
			5831: begin bcd3<=5;bcd2<=8;bcd1<=3;bcd0<=1; end
			5832: begin bcd3<=5;bcd2<=8;bcd1<=3;bcd0<=2; end
			5833: begin bcd3<=5;bcd2<=8;bcd1<=3;bcd0<=3; end
			5834: begin bcd3<=5;bcd2<=8;bcd1<=3;bcd0<=4; end
			5835: begin bcd3<=5;bcd2<=8;bcd1<=3;bcd0<=5; end
			5836: begin bcd3<=5;bcd2<=8;bcd1<=3;bcd0<=6; end
			5837: begin bcd3<=5;bcd2<=8;bcd1<=3;bcd0<=7; end
			5838: begin bcd3<=5;bcd2<=8;bcd1<=3;bcd0<=8; end
			5839: begin bcd3<=5;bcd2<=8;bcd1<=3;bcd0<=9; end
			5840: begin bcd3<=5;bcd2<=8;bcd1<=4;bcd0<=0; end
			5841: begin bcd3<=5;bcd2<=8;bcd1<=4;bcd0<=1; end
			5842: begin bcd3<=5;bcd2<=8;bcd1<=4;bcd0<=2; end
			5843: begin bcd3<=5;bcd2<=8;bcd1<=4;bcd0<=3; end
			5844: begin bcd3<=5;bcd2<=8;bcd1<=4;bcd0<=4; end
			5845: begin bcd3<=5;bcd2<=8;bcd1<=4;bcd0<=5; end
			5846: begin bcd3<=5;bcd2<=8;bcd1<=4;bcd0<=6; end
			5847: begin bcd3<=5;bcd2<=8;bcd1<=4;bcd0<=7; end
			5848: begin bcd3<=5;bcd2<=8;bcd1<=4;bcd0<=8; end
			5849: begin bcd3<=5;bcd2<=8;bcd1<=4;bcd0<=9; end
			5850: begin bcd3<=5;bcd2<=8;bcd1<=5;bcd0<=0; end
			5851: begin bcd3<=5;bcd2<=8;bcd1<=5;bcd0<=1; end
			5852: begin bcd3<=5;bcd2<=8;bcd1<=5;bcd0<=2; end
			5853: begin bcd3<=5;bcd2<=8;bcd1<=5;bcd0<=3; end
			5854: begin bcd3<=5;bcd2<=8;bcd1<=5;bcd0<=4; end
			5855: begin bcd3<=5;bcd2<=8;bcd1<=5;bcd0<=5; end
			5856: begin bcd3<=5;bcd2<=8;bcd1<=5;bcd0<=6; end
			5857: begin bcd3<=5;bcd2<=8;bcd1<=5;bcd0<=7; end
			5858: begin bcd3<=5;bcd2<=8;bcd1<=5;bcd0<=8; end
			5859: begin bcd3<=5;bcd2<=8;bcd1<=5;bcd0<=9; end
			5860: begin bcd3<=5;bcd2<=8;bcd1<=6;bcd0<=0; end
			5861: begin bcd3<=5;bcd2<=8;bcd1<=6;bcd0<=1; end
			5862: begin bcd3<=5;bcd2<=8;bcd1<=6;bcd0<=2; end
			5863: begin bcd3<=5;bcd2<=8;bcd1<=6;bcd0<=3; end
			5864: begin bcd3<=5;bcd2<=8;bcd1<=6;bcd0<=4; end
			5865: begin bcd3<=5;bcd2<=8;bcd1<=6;bcd0<=5; end
			5866: begin bcd3<=5;bcd2<=8;bcd1<=6;bcd0<=6; end
			5867: begin bcd3<=5;bcd2<=8;bcd1<=6;bcd0<=7; end
			5868: begin bcd3<=5;bcd2<=8;bcd1<=6;bcd0<=8; end
			5869: begin bcd3<=5;bcd2<=8;bcd1<=6;bcd0<=9; end
			5870: begin bcd3<=5;bcd2<=8;bcd1<=7;bcd0<=0; end
			5871: begin bcd3<=5;bcd2<=8;bcd1<=7;bcd0<=1; end
			5872: begin bcd3<=5;bcd2<=8;bcd1<=7;bcd0<=2; end
			5873: begin bcd3<=5;bcd2<=8;bcd1<=7;bcd0<=3; end
			5874: begin bcd3<=5;bcd2<=8;bcd1<=7;bcd0<=4; end
			5875: begin bcd3<=5;bcd2<=8;bcd1<=7;bcd0<=5; end
			5876: begin bcd3<=5;bcd2<=8;bcd1<=7;bcd0<=6; end
			5877: begin bcd3<=5;bcd2<=8;bcd1<=7;bcd0<=7; end
			5878: begin bcd3<=5;bcd2<=8;bcd1<=7;bcd0<=8; end
			5879: begin bcd3<=5;bcd2<=8;bcd1<=7;bcd0<=9; end
			5880: begin bcd3<=5;bcd2<=8;bcd1<=8;bcd0<=0; end
			5881: begin bcd3<=5;bcd2<=8;bcd1<=8;bcd0<=1; end
			5882: begin bcd3<=5;bcd2<=8;bcd1<=8;bcd0<=2; end
			5883: begin bcd3<=5;bcd2<=8;bcd1<=8;bcd0<=3; end
			5884: begin bcd3<=5;bcd2<=8;bcd1<=8;bcd0<=4; end
			5885: begin bcd3<=5;bcd2<=8;bcd1<=8;bcd0<=5; end
			5886: begin bcd3<=5;bcd2<=8;bcd1<=8;bcd0<=6; end
			5887: begin bcd3<=5;bcd2<=8;bcd1<=8;bcd0<=7; end
			5888: begin bcd3<=5;bcd2<=8;bcd1<=8;bcd0<=8; end
			5889: begin bcd3<=5;bcd2<=8;bcd1<=8;bcd0<=9; end
			5890: begin bcd3<=5;bcd2<=8;bcd1<=9;bcd0<=0; end
			5891: begin bcd3<=5;bcd2<=8;bcd1<=9;bcd0<=1; end
			5892: begin bcd3<=5;bcd2<=8;bcd1<=9;bcd0<=2; end
			5893: begin bcd3<=5;bcd2<=8;bcd1<=9;bcd0<=3; end
			5894: begin bcd3<=5;bcd2<=8;bcd1<=9;bcd0<=4; end
			5895: begin bcd3<=5;bcd2<=8;bcd1<=9;bcd0<=5; end
			5896: begin bcd3<=5;bcd2<=8;bcd1<=9;bcd0<=6; end
			5897: begin bcd3<=5;bcd2<=8;bcd1<=9;bcd0<=7; end
			5898: begin bcd3<=5;bcd2<=8;bcd1<=9;bcd0<=8; end
			5899: begin bcd3<=5;bcd2<=8;bcd1<=9;bcd0<=9; end
			5900: begin bcd3<=5;bcd2<=9;bcd1<=0;bcd0<=0; end
			5901: begin bcd3<=5;bcd2<=9;bcd1<=0;bcd0<=1; end
			5902: begin bcd3<=5;bcd2<=9;bcd1<=0;bcd0<=2; end
			5903: begin bcd3<=5;bcd2<=9;bcd1<=0;bcd0<=3; end
			5904: begin bcd3<=5;bcd2<=9;bcd1<=0;bcd0<=4; end
			5905: begin bcd3<=5;bcd2<=9;bcd1<=0;bcd0<=5; end
			5906: begin bcd3<=5;bcd2<=9;bcd1<=0;bcd0<=6; end
			5907: begin bcd3<=5;bcd2<=9;bcd1<=0;bcd0<=7; end
			5908: begin bcd3<=5;bcd2<=9;bcd1<=0;bcd0<=8; end
			5909: begin bcd3<=5;bcd2<=9;bcd1<=0;bcd0<=9; end
			5910: begin bcd3<=5;bcd2<=9;bcd1<=1;bcd0<=0; end
			5911: begin bcd3<=5;bcd2<=9;bcd1<=1;bcd0<=1; end
			5912: begin bcd3<=5;bcd2<=9;bcd1<=1;bcd0<=2; end
			5913: begin bcd3<=5;bcd2<=9;bcd1<=1;bcd0<=3; end
			5914: begin bcd3<=5;bcd2<=9;bcd1<=1;bcd0<=4; end
			5915: begin bcd3<=5;bcd2<=9;bcd1<=1;bcd0<=5; end
			5916: begin bcd3<=5;bcd2<=9;bcd1<=1;bcd0<=6; end
			5917: begin bcd3<=5;bcd2<=9;bcd1<=1;bcd0<=7; end
			5918: begin bcd3<=5;bcd2<=9;bcd1<=1;bcd0<=8; end
			5919: begin bcd3<=5;bcd2<=9;bcd1<=1;bcd0<=9; end
			5920: begin bcd3<=5;bcd2<=9;bcd1<=2;bcd0<=0; end
			5921: begin bcd3<=5;bcd2<=9;bcd1<=2;bcd0<=1; end
			5922: begin bcd3<=5;bcd2<=9;bcd1<=2;bcd0<=2; end
			5923: begin bcd3<=5;bcd2<=9;bcd1<=2;bcd0<=3; end
			5924: begin bcd3<=5;bcd2<=9;bcd1<=2;bcd0<=4; end
			5925: begin bcd3<=5;bcd2<=9;bcd1<=2;bcd0<=5; end
			5926: begin bcd3<=5;bcd2<=9;bcd1<=2;bcd0<=6; end
			5927: begin bcd3<=5;bcd2<=9;bcd1<=2;bcd0<=7; end
			5928: begin bcd3<=5;bcd2<=9;bcd1<=2;bcd0<=8; end
			5929: begin bcd3<=5;bcd2<=9;bcd1<=2;bcd0<=9; end
			5930: begin bcd3<=5;bcd2<=9;bcd1<=3;bcd0<=0; end
			5931: begin bcd3<=5;bcd2<=9;bcd1<=3;bcd0<=1; end
			5932: begin bcd3<=5;bcd2<=9;bcd1<=3;bcd0<=2; end
			5933: begin bcd3<=5;bcd2<=9;bcd1<=3;bcd0<=3; end
			5934: begin bcd3<=5;bcd2<=9;bcd1<=3;bcd0<=4; end
			5935: begin bcd3<=5;bcd2<=9;bcd1<=3;bcd0<=5; end
			5936: begin bcd3<=5;bcd2<=9;bcd1<=3;bcd0<=6; end
			5937: begin bcd3<=5;bcd2<=9;bcd1<=3;bcd0<=7; end
			5938: begin bcd3<=5;bcd2<=9;bcd1<=3;bcd0<=8; end
			5939: begin bcd3<=5;bcd2<=9;bcd1<=3;bcd0<=9; end
			5940: begin bcd3<=5;bcd2<=9;bcd1<=4;bcd0<=0; end
			5941: begin bcd3<=5;bcd2<=9;bcd1<=4;bcd0<=1; end
			5942: begin bcd3<=5;bcd2<=9;bcd1<=4;bcd0<=2; end
			5943: begin bcd3<=5;bcd2<=9;bcd1<=4;bcd0<=3; end
			5944: begin bcd3<=5;bcd2<=9;bcd1<=4;bcd0<=4; end
			5945: begin bcd3<=5;bcd2<=9;bcd1<=4;bcd0<=5; end
			5946: begin bcd3<=5;bcd2<=9;bcd1<=4;bcd0<=6; end
			5947: begin bcd3<=5;bcd2<=9;bcd1<=4;bcd0<=7; end
			5948: begin bcd3<=5;bcd2<=9;bcd1<=4;bcd0<=8; end
			5949: begin bcd3<=5;bcd2<=9;bcd1<=4;bcd0<=9; end
			5950: begin bcd3<=5;bcd2<=9;bcd1<=5;bcd0<=0; end
			5951: begin bcd3<=5;bcd2<=9;bcd1<=5;bcd0<=1; end
			5952: begin bcd3<=5;bcd2<=9;bcd1<=5;bcd0<=2; end
			5953: begin bcd3<=5;bcd2<=9;bcd1<=5;bcd0<=3; end
			5954: begin bcd3<=5;bcd2<=9;bcd1<=5;bcd0<=4; end
			5955: begin bcd3<=5;bcd2<=9;bcd1<=5;bcd0<=5; end
			5956: begin bcd3<=5;bcd2<=9;bcd1<=5;bcd0<=6; end
			5957: begin bcd3<=5;bcd2<=9;bcd1<=5;bcd0<=7; end
			5958: begin bcd3<=5;bcd2<=9;bcd1<=5;bcd0<=8; end
			5959: begin bcd3<=5;bcd2<=9;bcd1<=5;bcd0<=9; end
			5960: begin bcd3<=5;bcd2<=9;bcd1<=6;bcd0<=0; end
			5961: begin bcd3<=5;bcd2<=9;bcd1<=6;bcd0<=1; end
			5962: begin bcd3<=5;bcd2<=9;bcd1<=6;bcd0<=2; end
			5963: begin bcd3<=5;bcd2<=9;bcd1<=6;bcd0<=3; end
			5964: begin bcd3<=5;bcd2<=9;bcd1<=6;bcd0<=4; end
			5965: begin bcd3<=5;bcd2<=9;bcd1<=6;bcd0<=5; end
			5966: begin bcd3<=5;bcd2<=9;bcd1<=6;bcd0<=6; end
			5967: begin bcd3<=5;bcd2<=9;bcd1<=6;bcd0<=7; end
			5968: begin bcd3<=5;bcd2<=9;bcd1<=6;bcd0<=8; end
			5969: begin bcd3<=5;bcd2<=9;bcd1<=6;bcd0<=9; end
			5970: begin bcd3<=5;bcd2<=9;bcd1<=7;bcd0<=0; end
			5971: begin bcd3<=5;bcd2<=9;bcd1<=7;bcd0<=1; end
			5972: begin bcd3<=5;bcd2<=9;bcd1<=7;bcd0<=2; end
			5973: begin bcd3<=5;bcd2<=9;bcd1<=7;bcd0<=3; end
			5974: begin bcd3<=5;bcd2<=9;bcd1<=7;bcd0<=4; end
			5975: begin bcd3<=5;bcd2<=9;bcd1<=7;bcd0<=5; end
			5976: begin bcd3<=5;bcd2<=9;bcd1<=7;bcd0<=6; end
			5977: begin bcd3<=5;bcd2<=9;bcd1<=7;bcd0<=7; end
			5978: begin bcd3<=5;bcd2<=9;bcd1<=7;bcd0<=8; end
			5979: begin bcd3<=5;bcd2<=9;bcd1<=7;bcd0<=9; end
			5980: begin bcd3<=5;bcd2<=9;bcd1<=8;bcd0<=0; end
			5981: begin bcd3<=5;bcd2<=9;bcd1<=8;bcd0<=1; end
			5982: begin bcd3<=5;bcd2<=9;bcd1<=8;bcd0<=2; end
			5983: begin bcd3<=5;bcd2<=9;bcd1<=8;bcd0<=3; end
			5984: begin bcd3<=5;bcd2<=9;bcd1<=8;bcd0<=4; end
			5985: begin bcd3<=5;bcd2<=9;bcd1<=8;bcd0<=5; end
			5986: begin bcd3<=5;bcd2<=9;bcd1<=8;bcd0<=6; end
			5987: begin bcd3<=5;bcd2<=9;bcd1<=8;bcd0<=7; end
			5988: begin bcd3<=5;bcd2<=9;bcd1<=8;bcd0<=8; end
			5989: begin bcd3<=5;bcd2<=9;bcd1<=8;bcd0<=9; end
			5990: begin bcd3<=5;bcd2<=9;bcd1<=9;bcd0<=0; end
			5991: begin bcd3<=5;bcd2<=9;bcd1<=9;bcd0<=1; end
			5992: begin bcd3<=5;bcd2<=9;bcd1<=9;bcd0<=2; end
			5993: begin bcd3<=5;bcd2<=9;bcd1<=9;bcd0<=3; end
			5994: begin bcd3<=5;bcd2<=9;bcd1<=9;bcd0<=4; end
			5995: begin bcd3<=5;bcd2<=9;bcd1<=9;bcd0<=5; end
			5996: begin bcd3<=5;bcd2<=9;bcd1<=9;bcd0<=6; end
			5997: begin bcd3<=5;bcd2<=9;bcd1<=9;bcd0<=7; end
			5998: begin bcd3<=5;bcd2<=9;bcd1<=9;bcd0<=8; end
			5999: begin bcd3<=5;bcd2<=9;bcd1<=9;bcd0<=9; end
			6000: begin bcd3<=6;bcd2<=0;bcd1<=0;bcd0<=0; end
			6001: begin bcd3<=6;bcd2<=0;bcd1<=0;bcd0<=1; end
			6002: begin bcd3<=6;bcd2<=0;bcd1<=0;bcd0<=2; end
			6003: begin bcd3<=6;bcd2<=0;bcd1<=0;bcd0<=3; end
			6004: begin bcd3<=6;bcd2<=0;bcd1<=0;bcd0<=4; end
			6005: begin bcd3<=6;bcd2<=0;bcd1<=0;bcd0<=5; end
			6006: begin bcd3<=6;bcd2<=0;bcd1<=0;bcd0<=6; end
			6007: begin bcd3<=6;bcd2<=0;bcd1<=0;bcd0<=7; end
			6008: begin bcd3<=6;bcd2<=0;bcd1<=0;bcd0<=8; end
			6009: begin bcd3<=6;bcd2<=0;bcd1<=0;bcd0<=9; end
			6010: begin bcd3<=6;bcd2<=0;bcd1<=1;bcd0<=0; end
			6011: begin bcd3<=6;bcd2<=0;bcd1<=1;bcd0<=1; end
			6012: begin bcd3<=6;bcd2<=0;bcd1<=1;bcd0<=2; end
			6013: begin bcd3<=6;bcd2<=0;bcd1<=1;bcd0<=3; end
			6014: begin bcd3<=6;bcd2<=0;bcd1<=1;bcd0<=4; end
			6015: begin bcd3<=6;bcd2<=0;bcd1<=1;bcd0<=5; end
			6016: begin bcd3<=6;bcd2<=0;bcd1<=1;bcd0<=6; end
			6017: begin bcd3<=6;bcd2<=0;bcd1<=1;bcd0<=7; end
			6018: begin bcd3<=6;bcd2<=0;bcd1<=1;bcd0<=8; end
			6019: begin bcd3<=6;bcd2<=0;bcd1<=1;bcd0<=9; end
			6020: begin bcd3<=6;bcd2<=0;bcd1<=2;bcd0<=0; end
			6021: begin bcd3<=6;bcd2<=0;bcd1<=2;bcd0<=1; end
			6022: begin bcd3<=6;bcd2<=0;bcd1<=2;bcd0<=2; end
			6023: begin bcd3<=6;bcd2<=0;bcd1<=2;bcd0<=3; end
			6024: begin bcd3<=6;bcd2<=0;bcd1<=2;bcd0<=4; end
			6025: begin bcd3<=6;bcd2<=0;bcd1<=2;bcd0<=5; end
			6026: begin bcd3<=6;bcd2<=0;bcd1<=2;bcd0<=6; end
			6027: begin bcd3<=6;bcd2<=0;bcd1<=2;bcd0<=7; end
			6028: begin bcd3<=6;bcd2<=0;bcd1<=2;bcd0<=8; end
			6029: begin bcd3<=6;bcd2<=0;bcd1<=2;bcd0<=9; end
			6030: begin bcd3<=6;bcd2<=0;bcd1<=3;bcd0<=0; end
			6031: begin bcd3<=6;bcd2<=0;bcd1<=3;bcd0<=1; end
			6032: begin bcd3<=6;bcd2<=0;bcd1<=3;bcd0<=2; end
			6033: begin bcd3<=6;bcd2<=0;bcd1<=3;bcd0<=3; end
			6034: begin bcd3<=6;bcd2<=0;bcd1<=3;bcd0<=4; end
			6035: begin bcd3<=6;bcd2<=0;bcd1<=3;bcd0<=5; end
			6036: begin bcd3<=6;bcd2<=0;bcd1<=3;bcd0<=6; end
			6037: begin bcd3<=6;bcd2<=0;bcd1<=3;bcd0<=7; end
			6038: begin bcd3<=6;bcd2<=0;bcd1<=3;bcd0<=8; end
			6039: begin bcd3<=6;bcd2<=0;bcd1<=3;bcd0<=9; end
			6040: begin bcd3<=6;bcd2<=0;bcd1<=4;bcd0<=0; end
			6041: begin bcd3<=6;bcd2<=0;bcd1<=4;bcd0<=1; end
			6042: begin bcd3<=6;bcd2<=0;bcd1<=4;bcd0<=2; end
			6043: begin bcd3<=6;bcd2<=0;bcd1<=4;bcd0<=3; end
			6044: begin bcd3<=6;bcd2<=0;bcd1<=4;bcd0<=4; end
			6045: begin bcd3<=6;bcd2<=0;bcd1<=4;bcd0<=5; end
			6046: begin bcd3<=6;bcd2<=0;bcd1<=4;bcd0<=6; end
			6047: begin bcd3<=6;bcd2<=0;bcd1<=4;bcd0<=7; end
			6048: begin bcd3<=6;bcd2<=0;bcd1<=4;bcd0<=8; end
			6049: begin bcd3<=6;bcd2<=0;bcd1<=4;bcd0<=9; end
			6050: begin bcd3<=6;bcd2<=0;bcd1<=5;bcd0<=0; end
			6051: begin bcd3<=6;bcd2<=0;bcd1<=5;bcd0<=1; end
			6052: begin bcd3<=6;bcd2<=0;bcd1<=5;bcd0<=2; end
			6053: begin bcd3<=6;bcd2<=0;bcd1<=5;bcd0<=3; end
			6054: begin bcd3<=6;bcd2<=0;bcd1<=5;bcd0<=4; end
			6055: begin bcd3<=6;bcd2<=0;bcd1<=5;bcd0<=5; end
			6056: begin bcd3<=6;bcd2<=0;bcd1<=5;bcd0<=6; end
			6057: begin bcd3<=6;bcd2<=0;bcd1<=5;bcd0<=7; end
			6058: begin bcd3<=6;bcd2<=0;bcd1<=5;bcd0<=8; end
			6059: begin bcd3<=6;bcd2<=0;bcd1<=5;bcd0<=9; end
			6060: begin bcd3<=6;bcd2<=0;bcd1<=6;bcd0<=0; end
			6061: begin bcd3<=6;bcd2<=0;bcd1<=6;bcd0<=1; end
			6062: begin bcd3<=6;bcd2<=0;bcd1<=6;bcd0<=2; end
			6063: begin bcd3<=6;bcd2<=0;bcd1<=6;bcd0<=3; end
			6064: begin bcd3<=6;bcd2<=0;bcd1<=6;bcd0<=4; end
			6065: begin bcd3<=6;bcd2<=0;bcd1<=6;bcd0<=5; end
			6066: begin bcd3<=6;bcd2<=0;bcd1<=6;bcd0<=6; end
			6067: begin bcd3<=6;bcd2<=0;bcd1<=6;bcd0<=7; end
			6068: begin bcd3<=6;bcd2<=0;bcd1<=6;bcd0<=8; end
			6069: begin bcd3<=6;bcd2<=0;bcd1<=6;bcd0<=9; end
			6070: begin bcd3<=6;bcd2<=0;bcd1<=7;bcd0<=0; end
			6071: begin bcd3<=6;bcd2<=0;bcd1<=7;bcd0<=1; end
			6072: begin bcd3<=6;bcd2<=0;bcd1<=7;bcd0<=2; end
			6073: begin bcd3<=6;bcd2<=0;bcd1<=7;bcd0<=3; end
			6074: begin bcd3<=6;bcd2<=0;bcd1<=7;bcd0<=4; end
			6075: begin bcd3<=6;bcd2<=0;bcd1<=7;bcd0<=5; end
			6076: begin bcd3<=6;bcd2<=0;bcd1<=7;bcd0<=6; end
			6077: begin bcd3<=6;bcd2<=0;bcd1<=7;bcd0<=7; end
			6078: begin bcd3<=6;bcd2<=0;bcd1<=7;bcd0<=8; end
			6079: begin bcd3<=6;bcd2<=0;bcd1<=7;bcd0<=9; end
			6080: begin bcd3<=6;bcd2<=0;bcd1<=8;bcd0<=0; end
			6081: begin bcd3<=6;bcd2<=0;bcd1<=8;bcd0<=1; end
			6082: begin bcd3<=6;bcd2<=0;bcd1<=8;bcd0<=2; end
			6083: begin bcd3<=6;bcd2<=0;bcd1<=8;bcd0<=3; end
			6084: begin bcd3<=6;bcd2<=0;bcd1<=8;bcd0<=4; end
			6085: begin bcd3<=6;bcd2<=0;bcd1<=8;bcd0<=5; end
			6086: begin bcd3<=6;bcd2<=0;bcd1<=8;bcd0<=6; end
			6087: begin bcd3<=6;bcd2<=0;bcd1<=8;bcd0<=7; end
			6088: begin bcd3<=6;bcd2<=0;bcd1<=8;bcd0<=8; end
			6089: begin bcd3<=6;bcd2<=0;bcd1<=8;bcd0<=9; end
			6090: begin bcd3<=6;bcd2<=0;bcd1<=9;bcd0<=0; end
			6091: begin bcd3<=6;bcd2<=0;bcd1<=9;bcd0<=1; end
			6092: begin bcd3<=6;bcd2<=0;bcd1<=9;bcd0<=2; end
			6093: begin bcd3<=6;bcd2<=0;bcd1<=9;bcd0<=3; end
			6094: begin bcd3<=6;bcd2<=0;bcd1<=9;bcd0<=4; end
			6095: begin bcd3<=6;bcd2<=0;bcd1<=9;bcd0<=5; end
			6096: begin bcd3<=6;bcd2<=0;bcd1<=9;bcd0<=6; end
			6097: begin bcd3<=6;bcd2<=0;bcd1<=9;bcd0<=7; end
			6098: begin bcd3<=6;bcd2<=0;bcd1<=9;bcd0<=8; end
			6099: begin bcd3<=6;bcd2<=0;bcd1<=9;bcd0<=9; end
			6100: begin bcd3<=6;bcd2<=1;bcd1<=0;bcd0<=0; end
			6101: begin bcd3<=6;bcd2<=1;bcd1<=0;bcd0<=1; end
			6102: begin bcd3<=6;bcd2<=1;bcd1<=0;bcd0<=2; end
			6103: begin bcd3<=6;bcd2<=1;bcd1<=0;bcd0<=3; end
			6104: begin bcd3<=6;bcd2<=1;bcd1<=0;bcd0<=4; end
			6105: begin bcd3<=6;bcd2<=1;bcd1<=0;bcd0<=5; end
			6106: begin bcd3<=6;bcd2<=1;bcd1<=0;bcd0<=6; end
			6107: begin bcd3<=6;bcd2<=1;bcd1<=0;bcd0<=7; end
			6108: begin bcd3<=6;bcd2<=1;bcd1<=0;bcd0<=8; end
			6109: begin bcd3<=6;bcd2<=1;bcd1<=0;bcd0<=9; end
			6110: begin bcd3<=6;bcd2<=1;bcd1<=1;bcd0<=0; end
			6111: begin bcd3<=6;bcd2<=1;bcd1<=1;bcd0<=1; end
			6112: begin bcd3<=6;bcd2<=1;bcd1<=1;bcd0<=2; end
			6113: begin bcd3<=6;bcd2<=1;bcd1<=1;bcd0<=3; end
			6114: begin bcd3<=6;bcd2<=1;bcd1<=1;bcd0<=4; end
			6115: begin bcd3<=6;bcd2<=1;bcd1<=1;bcd0<=5; end
			6116: begin bcd3<=6;bcd2<=1;bcd1<=1;bcd0<=6; end
			6117: begin bcd3<=6;bcd2<=1;bcd1<=1;bcd0<=7; end
			6118: begin bcd3<=6;bcd2<=1;bcd1<=1;bcd0<=8; end
			6119: begin bcd3<=6;bcd2<=1;bcd1<=1;bcd0<=9; end
			6120: begin bcd3<=6;bcd2<=1;bcd1<=2;bcd0<=0; end
			6121: begin bcd3<=6;bcd2<=1;bcd1<=2;bcd0<=1; end
			6122: begin bcd3<=6;bcd2<=1;bcd1<=2;bcd0<=2; end
			6123: begin bcd3<=6;bcd2<=1;bcd1<=2;bcd0<=3; end
			6124: begin bcd3<=6;bcd2<=1;bcd1<=2;bcd0<=4; end
			6125: begin bcd3<=6;bcd2<=1;bcd1<=2;bcd0<=5; end
			6126: begin bcd3<=6;bcd2<=1;bcd1<=2;bcd0<=6; end
			6127: begin bcd3<=6;bcd2<=1;bcd1<=2;bcd0<=7; end
			6128: begin bcd3<=6;bcd2<=1;bcd1<=2;bcd0<=8; end
			6129: begin bcd3<=6;bcd2<=1;bcd1<=2;bcd0<=9; end
			6130: begin bcd3<=6;bcd2<=1;bcd1<=3;bcd0<=0; end
			6131: begin bcd3<=6;bcd2<=1;bcd1<=3;bcd0<=1; end
			6132: begin bcd3<=6;bcd2<=1;bcd1<=3;bcd0<=2; end
			6133: begin bcd3<=6;bcd2<=1;bcd1<=3;bcd0<=3; end
			6134: begin bcd3<=6;bcd2<=1;bcd1<=3;bcd0<=4; end
			6135: begin bcd3<=6;bcd2<=1;bcd1<=3;bcd0<=5; end
			6136: begin bcd3<=6;bcd2<=1;bcd1<=3;bcd0<=6; end
			6137: begin bcd3<=6;bcd2<=1;bcd1<=3;bcd0<=7; end
			6138: begin bcd3<=6;bcd2<=1;bcd1<=3;bcd0<=8; end
			6139: begin bcd3<=6;bcd2<=1;bcd1<=3;bcd0<=9; end
			6140: begin bcd3<=6;bcd2<=1;bcd1<=4;bcd0<=0; end
			6141: begin bcd3<=6;bcd2<=1;bcd1<=4;bcd0<=1; end
			6142: begin bcd3<=6;bcd2<=1;bcd1<=4;bcd0<=2; end
			6143: begin bcd3<=6;bcd2<=1;bcd1<=4;bcd0<=3; end
			6144: begin bcd3<=6;bcd2<=1;bcd1<=4;bcd0<=4; end
			6145: begin bcd3<=6;bcd2<=1;bcd1<=4;bcd0<=5; end
			6146: begin bcd3<=6;bcd2<=1;bcd1<=4;bcd0<=6; end
			6147: begin bcd3<=6;bcd2<=1;bcd1<=4;bcd0<=7; end
			6148: begin bcd3<=6;bcd2<=1;bcd1<=4;bcd0<=8; end
			6149: begin bcd3<=6;bcd2<=1;bcd1<=4;bcd0<=9; end
			6150: begin bcd3<=6;bcd2<=1;bcd1<=5;bcd0<=0; end
			6151: begin bcd3<=6;bcd2<=1;bcd1<=5;bcd0<=1; end
			6152: begin bcd3<=6;bcd2<=1;bcd1<=5;bcd0<=2; end
			6153: begin bcd3<=6;bcd2<=1;bcd1<=5;bcd0<=3; end
			6154: begin bcd3<=6;bcd2<=1;bcd1<=5;bcd0<=4; end
			6155: begin bcd3<=6;bcd2<=1;bcd1<=5;bcd0<=5; end
			6156: begin bcd3<=6;bcd2<=1;bcd1<=5;bcd0<=6; end
			6157: begin bcd3<=6;bcd2<=1;bcd1<=5;bcd0<=7; end
			6158: begin bcd3<=6;bcd2<=1;bcd1<=5;bcd0<=8; end
			6159: begin bcd3<=6;bcd2<=1;bcd1<=5;bcd0<=9; end
			6160: begin bcd3<=6;bcd2<=1;bcd1<=6;bcd0<=0; end
			6161: begin bcd3<=6;bcd2<=1;bcd1<=6;bcd0<=1; end
			6162: begin bcd3<=6;bcd2<=1;bcd1<=6;bcd0<=2; end
			6163: begin bcd3<=6;bcd2<=1;bcd1<=6;bcd0<=3; end
			6164: begin bcd3<=6;bcd2<=1;bcd1<=6;bcd0<=4; end
			6165: begin bcd3<=6;bcd2<=1;bcd1<=6;bcd0<=5; end
			6166: begin bcd3<=6;bcd2<=1;bcd1<=6;bcd0<=6; end
			6167: begin bcd3<=6;bcd2<=1;bcd1<=6;bcd0<=7; end
			6168: begin bcd3<=6;bcd2<=1;bcd1<=6;bcd0<=8; end
			6169: begin bcd3<=6;bcd2<=1;bcd1<=6;bcd0<=9; end
			6170: begin bcd3<=6;bcd2<=1;bcd1<=7;bcd0<=0; end
			6171: begin bcd3<=6;bcd2<=1;bcd1<=7;bcd0<=1; end
			6172: begin bcd3<=6;bcd2<=1;bcd1<=7;bcd0<=2; end
			6173: begin bcd3<=6;bcd2<=1;bcd1<=7;bcd0<=3; end
			6174: begin bcd3<=6;bcd2<=1;bcd1<=7;bcd0<=4; end
			6175: begin bcd3<=6;bcd2<=1;bcd1<=7;bcd0<=5; end
			6176: begin bcd3<=6;bcd2<=1;bcd1<=7;bcd0<=6; end
			6177: begin bcd3<=6;bcd2<=1;bcd1<=7;bcd0<=7; end
			6178: begin bcd3<=6;bcd2<=1;bcd1<=7;bcd0<=8; end
			6179: begin bcd3<=6;bcd2<=1;bcd1<=7;bcd0<=9; end
			6180: begin bcd3<=6;bcd2<=1;bcd1<=8;bcd0<=0; end
			6181: begin bcd3<=6;bcd2<=1;bcd1<=8;bcd0<=1; end
			6182: begin bcd3<=6;bcd2<=1;bcd1<=8;bcd0<=2; end
			6183: begin bcd3<=6;bcd2<=1;bcd1<=8;bcd0<=3; end
			6184: begin bcd3<=6;bcd2<=1;bcd1<=8;bcd0<=4; end
			6185: begin bcd3<=6;bcd2<=1;bcd1<=8;bcd0<=5; end
			6186: begin bcd3<=6;bcd2<=1;bcd1<=8;bcd0<=6; end
			6187: begin bcd3<=6;bcd2<=1;bcd1<=8;bcd0<=7; end
			6188: begin bcd3<=6;bcd2<=1;bcd1<=8;bcd0<=8; end
			6189: begin bcd3<=6;bcd2<=1;bcd1<=8;bcd0<=9; end
			6190: begin bcd3<=6;bcd2<=1;bcd1<=9;bcd0<=0; end
			6191: begin bcd3<=6;bcd2<=1;bcd1<=9;bcd0<=1; end
			6192: begin bcd3<=6;bcd2<=1;bcd1<=9;bcd0<=2; end
			6193: begin bcd3<=6;bcd2<=1;bcd1<=9;bcd0<=3; end
			6194: begin bcd3<=6;bcd2<=1;bcd1<=9;bcd0<=4; end
			6195: begin bcd3<=6;bcd2<=1;bcd1<=9;bcd0<=5; end
			6196: begin bcd3<=6;bcd2<=1;bcd1<=9;bcd0<=6; end
			6197: begin bcd3<=6;bcd2<=1;bcd1<=9;bcd0<=7; end
			6198: begin bcd3<=6;bcd2<=1;bcd1<=9;bcd0<=8; end
			6199: begin bcd3<=6;bcd2<=1;bcd1<=9;bcd0<=9; end
			6200: begin bcd3<=6;bcd2<=2;bcd1<=0;bcd0<=0; end
			6201: begin bcd3<=6;bcd2<=2;bcd1<=0;bcd0<=1; end
			6202: begin bcd3<=6;bcd2<=2;bcd1<=0;bcd0<=2; end
			6203: begin bcd3<=6;bcd2<=2;bcd1<=0;bcd0<=3; end
			6204: begin bcd3<=6;bcd2<=2;bcd1<=0;bcd0<=4; end
			6205: begin bcd3<=6;bcd2<=2;bcd1<=0;bcd0<=5; end
			6206: begin bcd3<=6;bcd2<=2;bcd1<=0;bcd0<=6; end
			6207: begin bcd3<=6;bcd2<=2;bcd1<=0;bcd0<=7; end
			6208: begin bcd3<=6;bcd2<=2;bcd1<=0;bcd0<=8; end
			6209: begin bcd3<=6;bcd2<=2;bcd1<=0;bcd0<=9; end
			6210: begin bcd3<=6;bcd2<=2;bcd1<=1;bcd0<=0; end
			6211: begin bcd3<=6;bcd2<=2;bcd1<=1;bcd0<=1; end
			6212: begin bcd3<=6;bcd2<=2;bcd1<=1;bcd0<=2; end
			6213: begin bcd3<=6;bcd2<=2;bcd1<=1;bcd0<=3; end
			6214: begin bcd3<=6;bcd2<=2;bcd1<=1;bcd0<=4; end
			6215: begin bcd3<=6;bcd2<=2;bcd1<=1;bcd0<=5; end
			6216: begin bcd3<=6;bcd2<=2;bcd1<=1;bcd0<=6; end
			6217: begin bcd3<=6;bcd2<=2;bcd1<=1;bcd0<=7; end
			6218: begin bcd3<=6;bcd2<=2;bcd1<=1;bcd0<=8; end
			6219: begin bcd3<=6;bcd2<=2;bcd1<=1;bcd0<=9; end
			6220: begin bcd3<=6;bcd2<=2;bcd1<=2;bcd0<=0; end
			6221: begin bcd3<=6;bcd2<=2;bcd1<=2;bcd0<=1; end
			6222: begin bcd3<=6;bcd2<=2;bcd1<=2;bcd0<=2; end
			6223: begin bcd3<=6;bcd2<=2;bcd1<=2;bcd0<=3; end
			6224: begin bcd3<=6;bcd2<=2;bcd1<=2;bcd0<=4; end
			6225: begin bcd3<=6;bcd2<=2;bcd1<=2;bcd0<=5; end
			6226: begin bcd3<=6;bcd2<=2;bcd1<=2;bcd0<=6; end
			6227: begin bcd3<=6;bcd2<=2;bcd1<=2;bcd0<=7; end
			6228: begin bcd3<=6;bcd2<=2;bcd1<=2;bcd0<=8; end
			6229: begin bcd3<=6;bcd2<=2;bcd1<=2;bcd0<=9; end
			6230: begin bcd3<=6;bcd2<=2;bcd1<=3;bcd0<=0; end
			6231: begin bcd3<=6;bcd2<=2;bcd1<=3;bcd0<=1; end
			6232: begin bcd3<=6;bcd2<=2;bcd1<=3;bcd0<=2; end
			6233: begin bcd3<=6;bcd2<=2;bcd1<=3;bcd0<=3; end
			6234: begin bcd3<=6;bcd2<=2;bcd1<=3;bcd0<=4; end
			6235: begin bcd3<=6;bcd2<=2;bcd1<=3;bcd0<=5; end
			6236: begin bcd3<=6;bcd2<=2;bcd1<=3;bcd0<=6; end
			6237: begin bcd3<=6;bcd2<=2;bcd1<=3;bcd0<=7; end
			6238: begin bcd3<=6;bcd2<=2;bcd1<=3;bcd0<=8; end
			6239: begin bcd3<=6;bcd2<=2;bcd1<=3;bcd0<=9; end
			6240: begin bcd3<=6;bcd2<=2;bcd1<=4;bcd0<=0; end
			6241: begin bcd3<=6;bcd2<=2;bcd1<=4;bcd0<=1; end
			6242: begin bcd3<=6;bcd2<=2;bcd1<=4;bcd0<=2; end
			6243: begin bcd3<=6;bcd2<=2;bcd1<=4;bcd0<=3; end
			6244: begin bcd3<=6;bcd2<=2;bcd1<=4;bcd0<=4; end
			6245: begin bcd3<=6;bcd2<=2;bcd1<=4;bcd0<=5; end
			6246: begin bcd3<=6;bcd2<=2;bcd1<=4;bcd0<=6; end
			6247: begin bcd3<=6;bcd2<=2;bcd1<=4;bcd0<=7; end
			6248: begin bcd3<=6;bcd2<=2;bcd1<=4;bcd0<=8; end
			6249: begin bcd3<=6;bcd2<=2;bcd1<=4;bcd0<=9; end
			6250: begin bcd3<=6;bcd2<=2;bcd1<=5;bcd0<=0; end
			6251: begin bcd3<=6;bcd2<=2;bcd1<=5;bcd0<=1; end
			6252: begin bcd3<=6;bcd2<=2;bcd1<=5;bcd0<=2; end
			6253: begin bcd3<=6;bcd2<=2;bcd1<=5;bcd0<=3; end
			6254: begin bcd3<=6;bcd2<=2;bcd1<=5;bcd0<=4; end
			6255: begin bcd3<=6;bcd2<=2;bcd1<=5;bcd0<=5; end
			6256: begin bcd3<=6;bcd2<=2;bcd1<=5;bcd0<=6; end
			6257: begin bcd3<=6;bcd2<=2;bcd1<=5;bcd0<=7; end
			6258: begin bcd3<=6;bcd2<=2;bcd1<=5;bcd0<=8; end
			6259: begin bcd3<=6;bcd2<=2;bcd1<=5;bcd0<=9; end
			6260: begin bcd3<=6;bcd2<=2;bcd1<=6;bcd0<=0; end
			6261: begin bcd3<=6;bcd2<=2;bcd1<=6;bcd0<=1; end
			6262: begin bcd3<=6;bcd2<=2;bcd1<=6;bcd0<=2; end
			6263: begin bcd3<=6;bcd2<=2;bcd1<=6;bcd0<=3; end
			6264: begin bcd3<=6;bcd2<=2;bcd1<=6;bcd0<=4; end
			6265: begin bcd3<=6;bcd2<=2;bcd1<=6;bcd0<=5; end
			6266: begin bcd3<=6;bcd2<=2;bcd1<=6;bcd0<=6; end
			6267: begin bcd3<=6;bcd2<=2;bcd1<=6;bcd0<=7; end
			6268: begin bcd3<=6;bcd2<=2;bcd1<=6;bcd0<=8; end
			6269: begin bcd3<=6;bcd2<=2;bcd1<=6;bcd0<=9; end
			6270: begin bcd3<=6;bcd2<=2;bcd1<=7;bcd0<=0; end
			6271: begin bcd3<=6;bcd2<=2;bcd1<=7;bcd0<=1; end
			6272: begin bcd3<=6;bcd2<=2;bcd1<=7;bcd0<=2; end
			6273: begin bcd3<=6;bcd2<=2;bcd1<=7;bcd0<=3; end
			6274: begin bcd3<=6;bcd2<=2;bcd1<=7;bcd0<=4; end
			6275: begin bcd3<=6;bcd2<=2;bcd1<=7;bcd0<=5; end
			6276: begin bcd3<=6;bcd2<=2;bcd1<=7;bcd0<=6; end
			6277: begin bcd3<=6;bcd2<=2;bcd1<=7;bcd0<=7; end
			6278: begin bcd3<=6;bcd2<=2;bcd1<=7;bcd0<=8; end
			6279: begin bcd3<=6;bcd2<=2;bcd1<=7;bcd0<=9; end
			6280: begin bcd3<=6;bcd2<=2;bcd1<=8;bcd0<=0; end
			6281: begin bcd3<=6;bcd2<=2;bcd1<=8;bcd0<=1; end
			6282: begin bcd3<=6;bcd2<=2;bcd1<=8;bcd0<=2; end
			6283: begin bcd3<=6;bcd2<=2;bcd1<=8;bcd0<=3; end
			6284: begin bcd3<=6;bcd2<=2;bcd1<=8;bcd0<=4; end
			6285: begin bcd3<=6;bcd2<=2;bcd1<=8;bcd0<=5; end
			6286: begin bcd3<=6;bcd2<=2;bcd1<=8;bcd0<=6; end
			6287: begin bcd3<=6;bcd2<=2;bcd1<=8;bcd0<=7; end
			6288: begin bcd3<=6;bcd2<=2;bcd1<=8;bcd0<=8; end
			6289: begin bcd3<=6;bcd2<=2;bcd1<=8;bcd0<=9; end
			6290: begin bcd3<=6;bcd2<=2;bcd1<=9;bcd0<=0; end
			6291: begin bcd3<=6;bcd2<=2;bcd1<=9;bcd0<=1; end
			6292: begin bcd3<=6;bcd2<=2;bcd1<=9;bcd0<=2; end
			6293: begin bcd3<=6;bcd2<=2;bcd1<=9;bcd0<=3; end
			6294: begin bcd3<=6;bcd2<=2;bcd1<=9;bcd0<=4; end
			6295: begin bcd3<=6;bcd2<=2;bcd1<=9;bcd0<=5; end
			6296: begin bcd3<=6;bcd2<=2;bcd1<=9;bcd0<=6; end
			6297: begin bcd3<=6;bcd2<=2;bcd1<=9;bcd0<=7; end
			6298: begin bcd3<=6;bcd2<=2;bcd1<=9;bcd0<=8; end
			6299: begin bcd3<=6;bcd2<=2;bcd1<=9;bcd0<=9; end
			6300: begin bcd3<=6;bcd2<=3;bcd1<=0;bcd0<=0; end
			6301: begin bcd3<=6;bcd2<=3;bcd1<=0;bcd0<=1; end
			6302: begin bcd3<=6;bcd2<=3;bcd1<=0;bcd0<=2; end
			6303: begin bcd3<=6;bcd2<=3;bcd1<=0;bcd0<=3; end
			6304: begin bcd3<=6;bcd2<=3;bcd1<=0;bcd0<=4; end
			6305: begin bcd3<=6;bcd2<=3;bcd1<=0;bcd0<=5; end
			6306: begin bcd3<=6;bcd2<=3;bcd1<=0;bcd0<=6; end
			6307: begin bcd3<=6;bcd2<=3;bcd1<=0;bcd0<=7; end
			6308: begin bcd3<=6;bcd2<=3;bcd1<=0;bcd0<=8; end
			6309: begin bcd3<=6;bcd2<=3;bcd1<=0;bcd0<=9; end
			6310: begin bcd3<=6;bcd2<=3;bcd1<=1;bcd0<=0; end
			6311: begin bcd3<=6;bcd2<=3;bcd1<=1;bcd0<=1; end
			6312: begin bcd3<=6;bcd2<=3;bcd1<=1;bcd0<=2; end
			6313: begin bcd3<=6;bcd2<=3;bcd1<=1;bcd0<=3; end
			6314: begin bcd3<=6;bcd2<=3;bcd1<=1;bcd0<=4; end
			6315: begin bcd3<=6;bcd2<=3;bcd1<=1;bcd0<=5; end
			6316: begin bcd3<=6;bcd2<=3;bcd1<=1;bcd0<=6; end
			6317: begin bcd3<=6;bcd2<=3;bcd1<=1;bcd0<=7; end
			6318: begin bcd3<=6;bcd2<=3;bcd1<=1;bcd0<=8; end
			6319: begin bcd3<=6;bcd2<=3;bcd1<=1;bcd0<=9; end
			6320: begin bcd3<=6;bcd2<=3;bcd1<=2;bcd0<=0; end
			6321: begin bcd3<=6;bcd2<=3;bcd1<=2;bcd0<=1; end
			6322: begin bcd3<=6;bcd2<=3;bcd1<=2;bcd0<=2; end
			6323: begin bcd3<=6;bcd2<=3;bcd1<=2;bcd0<=3; end
			6324: begin bcd3<=6;bcd2<=3;bcd1<=2;bcd0<=4; end
			6325: begin bcd3<=6;bcd2<=3;bcd1<=2;bcd0<=5; end
			6326: begin bcd3<=6;bcd2<=3;bcd1<=2;bcd0<=6; end
			6327: begin bcd3<=6;bcd2<=3;bcd1<=2;bcd0<=7; end
			6328: begin bcd3<=6;bcd2<=3;bcd1<=2;bcd0<=8; end
			6329: begin bcd3<=6;bcd2<=3;bcd1<=2;bcd0<=9; end
			6330: begin bcd3<=6;bcd2<=3;bcd1<=3;bcd0<=0; end
			6331: begin bcd3<=6;bcd2<=3;bcd1<=3;bcd0<=1; end
			6332: begin bcd3<=6;bcd2<=3;bcd1<=3;bcd0<=2; end
			6333: begin bcd3<=6;bcd2<=3;bcd1<=3;bcd0<=3; end
			6334: begin bcd3<=6;bcd2<=3;bcd1<=3;bcd0<=4; end
			6335: begin bcd3<=6;bcd2<=3;bcd1<=3;bcd0<=5; end
			6336: begin bcd3<=6;bcd2<=3;bcd1<=3;bcd0<=6; end
			6337: begin bcd3<=6;bcd2<=3;bcd1<=3;bcd0<=7; end
			6338: begin bcd3<=6;bcd2<=3;bcd1<=3;bcd0<=8; end
			6339: begin bcd3<=6;bcd2<=3;bcd1<=3;bcd0<=9; end
			6340: begin bcd3<=6;bcd2<=3;bcd1<=4;bcd0<=0; end
			6341: begin bcd3<=6;bcd2<=3;bcd1<=4;bcd0<=1; end
			6342: begin bcd3<=6;bcd2<=3;bcd1<=4;bcd0<=2; end
			6343: begin bcd3<=6;bcd2<=3;bcd1<=4;bcd0<=3; end
			6344: begin bcd3<=6;bcd2<=3;bcd1<=4;bcd0<=4; end
			6345: begin bcd3<=6;bcd2<=3;bcd1<=4;bcd0<=5; end
			6346: begin bcd3<=6;bcd2<=3;bcd1<=4;bcd0<=6; end
			6347: begin bcd3<=6;bcd2<=3;bcd1<=4;bcd0<=7; end
			6348: begin bcd3<=6;bcd2<=3;bcd1<=4;bcd0<=8; end
			6349: begin bcd3<=6;bcd2<=3;bcd1<=4;bcd0<=9; end
			6350: begin bcd3<=6;bcd2<=3;bcd1<=5;bcd0<=0; end
			6351: begin bcd3<=6;bcd2<=3;bcd1<=5;bcd0<=1; end
			6352: begin bcd3<=6;bcd2<=3;bcd1<=5;bcd0<=2; end
			6353: begin bcd3<=6;bcd2<=3;bcd1<=5;bcd0<=3; end
			6354: begin bcd3<=6;bcd2<=3;bcd1<=5;bcd0<=4; end
			6355: begin bcd3<=6;bcd2<=3;bcd1<=5;bcd0<=5; end
			6356: begin bcd3<=6;bcd2<=3;bcd1<=5;bcd0<=6; end
			6357: begin bcd3<=6;bcd2<=3;bcd1<=5;bcd0<=7; end
			6358: begin bcd3<=6;bcd2<=3;bcd1<=5;bcd0<=8; end
			6359: begin bcd3<=6;bcd2<=3;bcd1<=5;bcd0<=9; end
			6360: begin bcd3<=6;bcd2<=3;bcd1<=6;bcd0<=0; end
			6361: begin bcd3<=6;bcd2<=3;bcd1<=6;bcd0<=1; end
			6362: begin bcd3<=6;bcd2<=3;bcd1<=6;bcd0<=2; end
			6363: begin bcd3<=6;bcd2<=3;bcd1<=6;bcd0<=3; end
			6364: begin bcd3<=6;bcd2<=3;bcd1<=6;bcd0<=4; end
			6365: begin bcd3<=6;bcd2<=3;bcd1<=6;bcd0<=5; end
			6366: begin bcd3<=6;bcd2<=3;bcd1<=6;bcd0<=6; end
			6367: begin bcd3<=6;bcd2<=3;bcd1<=6;bcd0<=7; end
			6368: begin bcd3<=6;bcd2<=3;bcd1<=6;bcd0<=8; end
			6369: begin bcd3<=6;bcd2<=3;bcd1<=6;bcd0<=9; end
			6370: begin bcd3<=6;bcd2<=3;bcd1<=7;bcd0<=0; end
			6371: begin bcd3<=6;bcd2<=3;bcd1<=7;bcd0<=1; end
			6372: begin bcd3<=6;bcd2<=3;bcd1<=7;bcd0<=2; end
			6373: begin bcd3<=6;bcd2<=3;bcd1<=7;bcd0<=3; end
			6374: begin bcd3<=6;bcd2<=3;bcd1<=7;bcd0<=4; end
			6375: begin bcd3<=6;bcd2<=3;bcd1<=7;bcd0<=5; end
			6376: begin bcd3<=6;bcd2<=3;bcd1<=7;bcd0<=6; end
			6377: begin bcd3<=6;bcd2<=3;bcd1<=7;bcd0<=7; end
			6378: begin bcd3<=6;bcd2<=3;bcd1<=7;bcd0<=8; end
			6379: begin bcd3<=6;bcd2<=3;bcd1<=7;bcd0<=9; end
			6380: begin bcd3<=6;bcd2<=3;bcd1<=8;bcd0<=0; end
			6381: begin bcd3<=6;bcd2<=3;bcd1<=8;bcd0<=1; end
			6382: begin bcd3<=6;bcd2<=3;bcd1<=8;bcd0<=2; end
			6383: begin bcd3<=6;bcd2<=3;bcd1<=8;bcd0<=3; end
			6384: begin bcd3<=6;bcd2<=3;bcd1<=8;bcd0<=4; end
			6385: begin bcd3<=6;bcd2<=3;bcd1<=8;bcd0<=5; end
			6386: begin bcd3<=6;bcd2<=3;bcd1<=8;bcd0<=6; end
			6387: begin bcd3<=6;bcd2<=3;bcd1<=8;bcd0<=7; end
			6388: begin bcd3<=6;bcd2<=3;bcd1<=8;bcd0<=8; end
			6389: begin bcd3<=6;bcd2<=3;bcd1<=8;bcd0<=9; end
			6390: begin bcd3<=6;bcd2<=3;bcd1<=9;bcd0<=0; end
			6391: begin bcd3<=6;bcd2<=3;bcd1<=9;bcd0<=1; end
			6392: begin bcd3<=6;bcd2<=3;bcd1<=9;bcd0<=2; end
			6393: begin bcd3<=6;bcd2<=3;bcd1<=9;bcd0<=3; end
			6394: begin bcd3<=6;bcd2<=3;bcd1<=9;bcd0<=4; end
			6395: begin bcd3<=6;bcd2<=3;bcd1<=9;bcd0<=5; end
			6396: begin bcd3<=6;bcd2<=3;bcd1<=9;bcd0<=6; end
			6397: begin bcd3<=6;bcd2<=3;bcd1<=9;bcd0<=7; end
			6398: begin bcd3<=6;bcd2<=3;bcd1<=9;bcd0<=8; end
			6399: begin bcd3<=6;bcd2<=3;bcd1<=9;bcd0<=9; end
			6400: begin bcd3<=6;bcd2<=4;bcd1<=0;bcd0<=0; end
			6401: begin bcd3<=6;bcd2<=4;bcd1<=0;bcd0<=1; end
			6402: begin bcd3<=6;bcd2<=4;bcd1<=0;bcd0<=2; end
			6403: begin bcd3<=6;bcd2<=4;bcd1<=0;bcd0<=3; end
			6404: begin bcd3<=6;bcd2<=4;bcd1<=0;bcd0<=4; end
			6405: begin bcd3<=6;bcd2<=4;bcd1<=0;bcd0<=5; end
			6406: begin bcd3<=6;bcd2<=4;bcd1<=0;bcd0<=6; end
			6407: begin bcd3<=6;bcd2<=4;bcd1<=0;bcd0<=7; end
			6408: begin bcd3<=6;bcd2<=4;bcd1<=0;bcd0<=8; end
			6409: begin bcd3<=6;bcd2<=4;bcd1<=0;bcd0<=9; end
			6410: begin bcd3<=6;bcd2<=4;bcd1<=1;bcd0<=0; end
			6411: begin bcd3<=6;bcd2<=4;bcd1<=1;bcd0<=1; end
			6412: begin bcd3<=6;bcd2<=4;bcd1<=1;bcd0<=2; end
			6413: begin bcd3<=6;bcd2<=4;bcd1<=1;bcd0<=3; end
			6414: begin bcd3<=6;bcd2<=4;bcd1<=1;bcd0<=4; end
			6415: begin bcd3<=6;bcd2<=4;bcd1<=1;bcd0<=5; end
			6416: begin bcd3<=6;bcd2<=4;bcd1<=1;bcd0<=6; end
			6417: begin bcd3<=6;bcd2<=4;bcd1<=1;bcd0<=7; end
			6418: begin bcd3<=6;bcd2<=4;bcd1<=1;bcd0<=8; end
			6419: begin bcd3<=6;bcd2<=4;bcd1<=1;bcd0<=9; end
			6420: begin bcd3<=6;bcd2<=4;bcd1<=2;bcd0<=0; end
			6421: begin bcd3<=6;bcd2<=4;bcd1<=2;bcd0<=1; end
			6422: begin bcd3<=6;bcd2<=4;bcd1<=2;bcd0<=2; end
			6423: begin bcd3<=6;bcd2<=4;bcd1<=2;bcd0<=3; end
			6424: begin bcd3<=6;bcd2<=4;bcd1<=2;bcd0<=4; end
			6425: begin bcd3<=6;bcd2<=4;bcd1<=2;bcd0<=5; end
			6426: begin bcd3<=6;bcd2<=4;bcd1<=2;bcd0<=6; end
			6427: begin bcd3<=6;bcd2<=4;bcd1<=2;bcd0<=7; end
			6428: begin bcd3<=6;bcd2<=4;bcd1<=2;bcd0<=8; end
			6429: begin bcd3<=6;bcd2<=4;bcd1<=2;bcd0<=9; end
			6430: begin bcd3<=6;bcd2<=4;bcd1<=3;bcd0<=0; end
			6431: begin bcd3<=6;bcd2<=4;bcd1<=3;bcd0<=1; end
			6432: begin bcd3<=6;bcd2<=4;bcd1<=3;bcd0<=2; end
			6433: begin bcd3<=6;bcd2<=4;bcd1<=3;bcd0<=3; end
			6434: begin bcd3<=6;bcd2<=4;bcd1<=3;bcd0<=4; end
			6435: begin bcd3<=6;bcd2<=4;bcd1<=3;bcd0<=5; end
			6436: begin bcd3<=6;bcd2<=4;bcd1<=3;bcd0<=6; end
			6437: begin bcd3<=6;bcd2<=4;bcd1<=3;bcd0<=7; end
			6438: begin bcd3<=6;bcd2<=4;bcd1<=3;bcd0<=8; end
			6439: begin bcd3<=6;bcd2<=4;bcd1<=3;bcd0<=9; end
			6440: begin bcd3<=6;bcd2<=4;bcd1<=4;bcd0<=0; end
			6441: begin bcd3<=6;bcd2<=4;bcd1<=4;bcd0<=1; end
			6442: begin bcd3<=6;bcd2<=4;bcd1<=4;bcd0<=2; end
			6443: begin bcd3<=6;bcd2<=4;bcd1<=4;bcd0<=3; end
			6444: begin bcd3<=6;bcd2<=4;bcd1<=4;bcd0<=4; end
			6445: begin bcd3<=6;bcd2<=4;bcd1<=4;bcd0<=5; end
			6446: begin bcd3<=6;bcd2<=4;bcd1<=4;bcd0<=6; end
			6447: begin bcd3<=6;bcd2<=4;bcd1<=4;bcd0<=7; end
			6448: begin bcd3<=6;bcd2<=4;bcd1<=4;bcd0<=8; end
			6449: begin bcd3<=6;bcd2<=4;bcd1<=4;bcd0<=9; end
			6450: begin bcd3<=6;bcd2<=4;bcd1<=5;bcd0<=0; end
			6451: begin bcd3<=6;bcd2<=4;bcd1<=5;bcd0<=1; end
			6452: begin bcd3<=6;bcd2<=4;bcd1<=5;bcd0<=2; end
			6453: begin bcd3<=6;bcd2<=4;bcd1<=5;bcd0<=3; end
			6454: begin bcd3<=6;bcd2<=4;bcd1<=5;bcd0<=4; end
			6455: begin bcd3<=6;bcd2<=4;bcd1<=5;bcd0<=5; end
			6456: begin bcd3<=6;bcd2<=4;bcd1<=5;bcd0<=6; end
			6457: begin bcd3<=6;bcd2<=4;bcd1<=5;bcd0<=7; end
			6458: begin bcd3<=6;bcd2<=4;bcd1<=5;bcd0<=8; end
			6459: begin bcd3<=6;bcd2<=4;bcd1<=5;bcd0<=9; end
			6460: begin bcd3<=6;bcd2<=4;bcd1<=6;bcd0<=0; end
			6461: begin bcd3<=6;bcd2<=4;bcd1<=6;bcd0<=1; end
			6462: begin bcd3<=6;bcd2<=4;bcd1<=6;bcd0<=2; end
			6463: begin bcd3<=6;bcd2<=4;bcd1<=6;bcd0<=3; end
			6464: begin bcd3<=6;bcd2<=4;bcd1<=6;bcd0<=4; end
			6465: begin bcd3<=6;bcd2<=4;bcd1<=6;bcd0<=5; end
			6466: begin bcd3<=6;bcd2<=4;bcd1<=6;bcd0<=6; end
			6467: begin bcd3<=6;bcd2<=4;bcd1<=6;bcd0<=7; end
			6468: begin bcd3<=6;bcd2<=4;bcd1<=6;bcd0<=8; end
			6469: begin bcd3<=6;bcd2<=4;bcd1<=6;bcd0<=9; end
			6470: begin bcd3<=6;bcd2<=4;bcd1<=7;bcd0<=0; end
			6471: begin bcd3<=6;bcd2<=4;bcd1<=7;bcd0<=1; end
			6472: begin bcd3<=6;bcd2<=4;bcd1<=7;bcd0<=2; end
			6473: begin bcd3<=6;bcd2<=4;bcd1<=7;bcd0<=3; end
			6474: begin bcd3<=6;bcd2<=4;bcd1<=7;bcd0<=4; end
			6475: begin bcd3<=6;bcd2<=4;bcd1<=7;bcd0<=5; end
			6476: begin bcd3<=6;bcd2<=4;bcd1<=7;bcd0<=6; end
			6477: begin bcd3<=6;bcd2<=4;bcd1<=7;bcd0<=7; end
			6478: begin bcd3<=6;bcd2<=4;bcd1<=7;bcd0<=8; end
			6479: begin bcd3<=6;bcd2<=4;bcd1<=7;bcd0<=9; end
			6480: begin bcd3<=6;bcd2<=4;bcd1<=8;bcd0<=0; end
			6481: begin bcd3<=6;bcd2<=4;bcd1<=8;bcd0<=1; end
			6482: begin bcd3<=6;bcd2<=4;bcd1<=8;bcd0<=2; end
			6483: begin bcd3<=6;bcd2<=4;bcd1<=8;bcd0<=3; end
			6484: begin bcd3<=6;bcd2<=4;bcd1<=8;bcd0<=4; end
			6485: begin bcd3<=6;bcd2<=4;bcd1<=8;bcd0<=5; end
			6486: begin bcd3<=6;bcd2<=4;bcd1<=8;bcd0<=6; end
			6487: begin bcd3<=6;bcd2<=4;bcd1<=8;bcd0<=7; end
			6488: begin bcd3<=6;bcd2<=4;bcd1<=8;bcd0<=8; end
			6489: begin bcd3<=6;bcd2<=4;bcd1<=8;bcd0<=9; end
			6490: begin bcd3<=6;bcd2<=4;bcd1<=9;bcd0<=0; end
			6491: begin bcd3<=6;bcd2<=4;bcd1<=9;bcd0<=1; end
			6492: begin bcd3<=6;bcd2<=4;bcd1<=9;bcd0<=2; end
			6493: begin bcd3<=6;bcd2<=4;bcd1<=9;bcd0<=3; end
			6494: begin bcd3<=6;bcd2<=4;bcd1<=9;bcd0<=4; end
			6495: begin bcd3<=6;bcd2<=4;bcd1<=9;bcd0<=5; end
			6496: begin bcd3<=6;bcd2<=4;bcd1<=9;bcd0<=6; end
			6497: begin bcd3<=6;bcd2<=4;bcd1<=9;bcd0<=7; end
			6498: begin bcd3<=6;bcd2<=4;bcd1<=9;bcd0<=8; end
			6499: begin bcd3<=6;bcd2<=4;bcd1<=9;bcd0<=9; end
			6500: begin bcd3<=6;bcd2<=5;bcd1<=0;bcd0<=0; end
			6501: begin bcd3<=6;bcd2<=5;bcd1<=0;bcd0<=1; end
			6502: begin bcd3<=6;bcd2<=5;bcd1<=0;bcd0<=2; end
			6503: begin bcd3<=6;bcd2<=5;bcd1<=0;bcd0<=3; end
			6504: begin bcd3<=6;bcd2<=5;bcd1<=0;bcd0<=4; end
			6505: begin bcd3<=6;bcd2<=5;bcd1<=0;bcd0<=5; end
			6506: begin bcd3<=6;bcd2<=5;bcd1<=0;bcd0<=6; end
			6507: begin bcd3<=6;bcd2<=5;bcd1<=0;bcd0<=7; end
			6508: begin bcd3<=6;bcd2<=5;bcd1<=0;bcd0<=8; end
			6509: begin bcd3<=6;bcd2<=5;bcd1<=0;bcd0<=9; end
			6510: begin bcd3<=6;bcd2<=5;bcd1<=1;bcd0<=0; end
			6511: begin bcd3<=6;bcd2<=5;bcd1<=1;bcd0<=1; end
			6512: begin bcd3<=6;bcd2<=5;bcd1<=1;bcd0<=2; end
			6513: begin bcd3<=6;bcd2<=5;bcd1<=1;bcd0<=3; end
			6514: begin bcd3<=6;bcd2<=5;bcd1<=1;bcd0<=4; end
			6515: begin bcd3<=6;bcd2<=5;bcd1<=1;bcd0<=5; end
			6516: begin bcd3<=6;bcd2<=5;bcd1<=1;bcd0<=6; end
			6517: begin bcd3<=6;bcd2<=5;bcd1<=1;bcd0<=7; end
			6518: begin bcd3<=6;bcd2<=5;bcd1<=1;bcd0<=8; end
			6519: begin bcd3<=6;bcd2<=5;bcd1<=1;bcd0<=9; end
			6520: begin bcd3<=6;bcd2<=5;bcd1<=2;bcd0<=0; end
			6521: begin bcd3<=6;bcd2<=5;bcd1<=2;bcd0<=1; end
			6522: begin bcd3<=6;bcd2<=5;bcd1<=2;bcd0<=2; end
			6523: begin bcd3<=6;bcd2<=5;bcd1<=2;bcd0<=3; end
			6524: begin bcd3<=6;bcd2<=5;bcd1<=2;bcd0<=4; end
			6525: begin bcd3<=6;bcd2<=5;bcd1<=2;bcd0<=5; end
			6526: begin bcd3<=6;bcd2<=5;bcd1<=2;bcd0<=6; end
			6527: begin bcd3<=6;bcd2<=5;bcd1<=2;bcd0<=7; end
			6528: begin bcd3<=6;bcd2<=5;bcd1<=2;bcd0<=8; end
			6529: begin bcd3<=6;bcd2<=5;bcd1<=2;bcd0<=9; end
			6530: begin bcd3<=6;bcd2<=5;bcd1<=3;bcd0<=0; end
			6531: begin bcd3<=6;bcd2<=5;bcd1<=3;bcd0<=1; end
			6532: begin bcd3<=6;bcd2<=5;bcd1<=3;bcd0<=2; end
			6533: begin bcd3<=6;bcd2<=5;bcd1<=3;bcd0<=3; end
			6534: begin bcd3<=6;bcd2<=5;bcd1<=3;bcd0<=4; end
			6535: begin bcd3<=6;bcd2<=5;bcd1<=3;bcd0<=5; end
			6536: begin bcd3<=6;bcd2<=5;bcd1<=3;bcd0<=6; end
			6537: begin bcd3<=6;bcd2<=5;bcd1<=3;bcd0<=7; end
			6538: begin bcd3<=6;bcd2<=5;bcd1<=3;bcd0<=8; end
			6539: begin bcd3<=6;bcd2<=5;bcd1<=3;bcd0<=9; end
			6540: begin bcd3<=6;bcd2<=5;bcd1<=4;bcd0<=0; end
			6541: begin bcd3<=6;bcd2<=5;bcd1<=4;bcd0<=1; end
			6542: begin bcd3<=6;bcd2<=5;bcd1<=4;bcd0<=2; end
			6543: begin bcd3<=6;bcd2<=5;bcd1<=4;bcd0<=3; end
			6544: begin bcd3<=6;bcd2<=5;bcd1<=4;bcd0<=4; end
			6545: begin bcd3<=6;bcd2<=5;bcd1<=4;bcd0<=5; end
			6546: begin bcd3<=6;bcd2<=5;bcd1<=4;bcd0<=6; end
			6547: begin bcd3<=6;bcd2<=5;bcd1<=4;bcd0<=7; end
			6548: begin bcd3<=6;bcd2<=5;bcd1<=4;bcd0<=8; end
			6549: begin bcd3<=6;bcd2<=5;bcd1<=4;bcd0<=9; end
			6550: begin bcd3<=6;bcd2<=5;bcd1<=5;bcd0<=0; end
			6551: begin bcd3<=6;bcd2<=5;bcd1<=5;bcd0<=1; end
			6552: begin bcd3<=6;bcd2<=5;bcd1<=5;bcd0<=2; end
			6553: begin bcd3<=6;bcd2<=5;bcd1<=5;bcd0<=3; end
			6554: begin bcd3<=6;bcd2<=5;bcd1<=5;bcd0<=4; end
			6555: begin bcd3<=6;bcd2<=5;bcd1<=5;bcd0<=5; end
			6556: begin bcd3<=6;bcd2<=5;bcd1<=5;bcd0<=6; end
			6557: begin bcd3<=6;bcd2<=5;bcd1<=5;bcd0<=7; end
			6558: begin bcd3<=6;bcd2<=5;bcd1<=5;bcd0<=8; end
			6559: begin bcd3<=6;bcd2<=5;bcd1<=5;bcd0<=9; end
			6560: begin bcd3<=6;bcd2<=5;bcd1<=6;bcd0<=0; end
			6561: begin bcd3<=6;bcd2<=5;bcd1<=6;bcd0<=1; end
			6562: begin bcd3<=6;bcd2<=5;bcd1<=6;bcd0<=2; end
			6563: begin bcd3<=6;bcd2<=5;bcd1<=6;bcd0<=3; end
			6564: begin bcd3<=6;bcd2<=5;bcd1<=6;bcd0<=4; end
			6565: begin bcd3<=6;bcd2<=5;bcd1<=6;bcd0<=5; end
			6566: begin bcd3<=6;bcd2<=5;bcd1<=6;bcd0<=6; end
			6567: begin bcd3<=6;bcd2<=5;bcd1<=6;bcd0<=7; end
			6568: begin bcd3<=6;bcd2<=5;bcd1<=6;bcd0<=8; end
			6569: begin bcd3<=6;bcd2<=5;bcd1<=6;bcd0<=9; end
			6570: begin bcd3<=6;bcd2<=5;bcd1<=7;bcd0<=0; end
			6571: begin bcd3<=6;bcd2<=5;bcd1<=7;bcd0<=1; end
			6572: begin bcd3<=6;bcd2<=5;bcd1<=7;bcd0<=2; end
			6573: begin bcd3<=6;bcd2<=5;bcd1<=7;bcd0<=3; end
			6574: begin bcd3<=6;bcd2<=5;bcd1<=7;bcd0<=4; end
			6575: begin bcd3<=6;bcd2<=5;bcd1<=7;bcd0<=5; end
			6576: begin bcd3<=6;bcd2<=5;bcd1<=7;bcd0<=6; end
			6577: begin bcd3<=6;bcd2<=5;bcd1<=7;bcd0<=7; end
			6578: begin bcd3<=6;bcd2<=5;bcd1<=7;bcd0<=8; end
			6579: begin bcd3<=6;bcd2<=5;bcd1<=7;bcd0<=9; end
			6580: begin bcd3<=6;bcd2<=5;bcd1<=8;bcd0<=0; end
			6581: begin bcd3<=6;bcd2<=5;bcd1<=8;bcd0<=1; end
			6582: begin bcd3<=6;bcd2<=5;bcd1<=8;bcd0<=2; end
			6583: begin bcd3<=6;bcd2<=5;bcd1<=8;bcd0<=3; end
			6584: begin bcd3<=6;bcd2<=5;bcd1<=8;bcd0<=4; end
			6585: begin bcd3<=6;bcd2<=5;bcd1<=8;bcd0<=5; end
			6586: begin bcd3<=6;bcd2<=5;bcd1<=8;bcd0<=6; end
			6587: begin bcd3<=6;bcd2<=5;bcd1<=8;bcd0<=7; end
			6588: begin bcd3<=6;bcd2<=5;bcd1<=8;bcd0<=8; end
			6589: begin bcd3<=6;bcd2<=5;bcd1<=8;bcd0<=9; end
			6590: begin bcd3<=6;bcd2<=5;bcd1<=9;bcd0<=0; end
			6591: begin bcd3<=6;bcd2<=5;bcd1<=9;bcd0<=1; end
			6592: begin bcd3<=6;bcd2<=5;bcd1<=9;bcd0<=2; end
			6593: begin bcd3<=6;bcd2<=5;bcd1<=9;bcd0<=3; end
			6594: begin bcd3<=6;bcd2<=5;bcd1<=9;bcd0<=4; end
			6595: begin bcd3<=6;bcd2<=5;bcd1<=9;bcd0<=5; end
			6596: begin bcd3<=6;bcd2<=5;bcd1<=9;bcd0<=6; end
			6597: begin bcd3<=6;bcd2<=5;bcd1<=9;bcd0<=7; end
			6598: begin bcd3<=6;bcd2<=5;bcd1<=9;bcd0<=8; end
			6599: begin bcd3<=6;bcd2<=5;bcd1<=9;bcd0<=9; end
			6600: begin bcd3<=6;bcd2<=6;bcd1<=0;bcd0<=0; end
			6601: begin bcd3<=6;bcd2<=6;bcd1<=0;bcd0<=1; end
			6602: begin bcd3<=6;bcd2<=6;bcd1<=0;bcd0<=2; end
			6603: begin bcd3<=6;bcd2<=6;bcd1<=0;bcd0<=3; end
			6604: begin bcd3<=6;bcd2<=6;bcd1<=0;bcd0<=4; end
			6605: begin bcd3<=6;bcd2<=6;bcd1<=0;bcd0<=5; end
			6606: begin bcd3<=6;bcd2<=6;bcd1<=0;bcd0<=6; end
			6607: begin bcd3<=6;bcd2<=6;bcd1<=0;bcd0<=7; end
			6608: begin bcd3<=6;bcd2<=6;bcd1<=0;bcd0<=8; end
			6609: begin bcd3<=6;bcd2<=6;bcd1<=0;bcd0<=9; end
			6610: begin bcd3<=6;bcd2<=6;bcd1<=1;bcd0<=0; end
			6611: begin bcd3<=6;bcd2<=6;bcd1<=1;bcd0<=1; end
			6612: begin bcd3<=6;bcd2<=6;bcd1<=1;bcd0<=2; end
			6613: begin bcd3<=6;bcd2<=6;bcd1<=1;bcd0<=3; end
			6614: begin bcd3<=6;bcd2<=6;bcd1<=1;bcd0<=4; end
			6615: begin bcd3<=6;bcd2<=6;bcd1<=1;bcd0<=5; end
			6616: begin bcd3<=6;bcd2<=6;bcd1<=1;bcd0<=6; end
			6617: begin bcd3<=6;bcd2<=6;bcd1<=1;bcd0<=7; end
			6618: begin bcd3<=6;bcd2<=6;bcd1<=1;bcd0<=8; end
			6619: begin bcd3<=6;bcd2<=6;bcd1<=1;bcd0<=9; end
			6620: begin bcd3<=6;bcd2<=6;bcd1<=2;bcd0<=0; end
			6621: begin bcd3<=6;bcd2<=6;bcd1<=2;bcd0<=1; end
			6622: begin bcd3<=6;bcd2<=6;bcd1<=2;bcd0<=2; end
			6623: begin bcd3<=6;bcd2<=6;bcd1<=2;bcd0<=3; end
			6624: begin bcd3<=6;bcd2<=6;bcd1<=2;bcd0<=4; end
			6625: begin bcd3<=6;bcd2<=6;bcd1<=2;bcd0<=5; end
			6626: begin bcd3<=6;bcd2<=6;bcd1<=2;bcd0<=6; end
			6627: begin bcd3<=6;bcd2<=6;bcd1<=2;bcd0<=7; end
			6628: begin bcd3<=6;bcd2<=6;bcd1<=2;bcd0<=8; end
			6629: begin bcd3<=6;bcd2<=6;bcd1<=2;bcd0<=9; end
			6630: begin bcd3<=6;bcd2<=6;bcd1<=3;bcd0<=0; end
			6631: begin bcd3<=6;bcd2<=6;bcd1<=3;bcd0<=1; end
			6632: begin bcd3<=6;bcd2<=6;bcd1<=3;bcd0<=2; end
			6633: begin bcd3<=6;bcd2<=6;bcd1<=3;bcd0<=3; end
			6634: begin bcd3<=6;bcd2<=6;bcd1<=3;bcd0<=4; end
			6635: begin bcd3<=6;bcd2<=6;bcd1<=3;bcd0<=5; end
			6636: begin bcd3<=6;bcd2<=6;bcd1<=3;bcd0<=6; end
			6637: begin bcd3<=6;bcd2<=6;bcd1<=3;bcd0<=7; end
			6638: begin bcd3<=6;bcd2<=6;bcd1<=3;bcd0<=8; end
			6639: begin bcd3<=6;bcd2<=6;bcd1<=3;bcd0<=9; end
			6640: begin bcd3<=6;bcd2<=6;bcd1<=4;bcd0<=0; end
			6641: begin bcd3<=6;bcd2<=6;bcd1<=4;bcd0<=1; end
			6642: begin bcd3<=6;bcd2<=6;bcd1<=4;bcd0<=2; end
			6643: begin bcd3<=6;bcd2<=6;bcd1<=4;bcd0<=3; end
			6644: begin bcd3<=6;bcd2<=6;bcd1<=4;bcd0<=4; end
			6645: begin bcd3<=6;bcd2<=6;bcd1<=4;bcd0<=5; end
			6646: begin bcd3<=6;bcd2<=6;bcd1<=4;bcd0<=6; end
			6647: begin bcd3<=6;bcd2<=6;bcd1<=4;bcd0<=7; end
			6648: begin bcd3<=6;bcd2<=6;bcd1<=4;bcd0<=8; end
			6649: begin bcd3<=6;bcd2<=6;bcd1<=4;bcd0<=9; end
			6650: begin bcd3<=6;bcd2<=6;bcd1<=5;bcd0<=0; end
			6651: begin bcd3<=6;bcd2<=6;bcd1<=5;bcd0<=1; end
			6652: begin bcd3<=6;bcd2<=6;bcd1<=5;bcd0<=2; end
			6653: begin bcd3<=6;bcd2<=6;bcd1<=5;bcd0<=3; end
			6654: begin bcd3<=6;bcd2<=6;bcd1<=5;bcd0<=4; end
			6655: begin bcd3<=6;bcd2<=6;bcd1<=5;bcd0<=5; end
			6656: begin bcd3<=6;bcd2<=6;bcd1<=5;bcd0<=6; end
			6657: begin bcd3<=6;bcd2<=6;bcd1<=5;bcd0<=7; end
			6658: begin bcd3<=6;bcd2<=6;bcd1<=5;bcd0<=8; end
			6659: begin bcd3<=6;bcd2<=6;bcd1<=5;bcd0<=9; end
			6660: begin bcd3<=6;bcd2<=6;bcd1<=6;bcd0<=0; end
			6661: begin bcd3<=6;bcd2<=6;bcd1<=6;bcd0<=1; end
			6662: begin bcd3<=6;bcd2<=6;bcd1<=6;bcd0<=2; end
			6663: begin bcd3<=6;bcd2<=6;bcd1<=6;bcd0<=3; end
			6664: begin bcd3<=6;bcd2<=6;bcd1<=6;bcd0<=4; end
			6665: begin bcd3<=6;bcd2<=6;bcd1<=6;bcd0<=5; end
			6666: begin bcd3<=6;bcd2<=6;bcd1<=6;bcd0<=6; end
			6667: begin bcd3<=6;bcd2<=6;bcd1<=6;bcd0<=7; end
			6668: begin bcd3<=6;bcd2<=6;bcd1<=6;bcd0<=8; end
			6669: begin bcd3<=6;bcd2<=6;bcd1<=6;bcd0<=9; end
			6670: begin bcd3<=6;bcd2<=6;bcd1<=7;bcd0<=0; end
			6671: begin bcd3<=6;bcd2<=6;bcd1<=7;bcd0<=1; end
			6672: begin bcd3<=6;bcd2<=6;bcd1<=7;bcd0<=2; end
			6673: begin bcd3<=6;bcd2<=6;bcd1<=7;bcd0<=3; end
			6674: begin bcd3<=6;bcd2<=6;bcd1<=7;bcd0<=4; end
			6675: begin bcd3<=6;bcd2<=6;bcd1<=7;bcd0<=5; end
			6676: begin bcd3<=6;bcd2<=6;bcd1<=7;bcd0<=6; end
			6677: begin bcd3<=6;bcd2<=6;bcd1<=7;bcd0<=7; end
			6678: begin bcd3<=6;bcd2<=6;bcd1<=7;bcd0<=8; end
			6679: begin bcd3<=6;bcd2<=6;bcd1<=7;bcd0<=9; end
			6680: begin bcd3<=6;bcd2<=6;bcd1<=8;bcd0<=0; end
			6681: begin bcd3<=6;bcd2<=6;bcd1<=8;bcd0<=1; end
			6682: begin bcd3<=6;bcd2<=6;bcd1<=8;bcd0<=2; end
			6683: begin bcd3<=6;bcd2<=6;bcd1<=8;bcd0<=3; end
			6684: begin bcd3<=6;bcd2<=6;bcd1<=8;bcd0<=4; end
			6685: begin bcd3<=6;bcd2<=6;bcd1<=8;bcd0<=5; end
			6686: begin bcd3<=6;bcd2<=6;bcd1<=8;bcd0<=6; end
			6687: begin bcd3<=6;bcd2<=6;bcd1<=8;bcd0<=7; end
			6688: begin bcd3<=6;bcd2<=6;bcd1<=8;bcd0<=8; end
			6689: begin bcd3<=6;bcd2<=6;bcd1<=8;bcd0<=9; end
			6690: begin bcd3<=6;bcd2<=6;bcd1<=9;bcd0<=0; end
			6691: begin bcd3<=6;bcd2<=6;bcd1<=9;bcd0<=1; end
			6692: begin bcd3<=6;bcd2<=6;bcd1<=9;bcd0<=2; end
			6693: begin bcd3<=6;bcd2<=6;bcd1<=9;bcd0<=3; end
			6694: begin bcd3<=6;bcd2<=6;bcd1<=9;bcd0<=4; end
			6695: begin bcd3<=6;bcd2<=6;bcd1<=9;bcd0<=5; end
			6696: begin bcd3<=6;bcd2<=6;bcd1<=9;bcd0<=6; end
			6697: begin bcd3<=6;bcd2<=6;bcd1<=9;bcd0<=7; end
			6698: begin bcd3<=6;bcd2<=6;bcd1<=9;bcd0<=8; end
			6699: begin bcd3<=6;bcd2<=6;bcd1<=9;bcd0<=9; end
			6700: begin bcd3<=6;bcd2<=7;bcd1<=0;bcd0<=0; end
			6701: begin bcd3<=6;bcd2<=7;bcd1<=0;bcd0<=1; end
			6702: begin bcd3<=6;bcd2<=7;bcd1<=0;bcd0<=2; end
			6703: begin bcd3<=6;bcd2<=7;bcd1<=0;bcd0<=3; end
			6704: begin bcd3<=6;bcd2<=7;bcd1<=0;bcd0<=4; end
			6705: begin bcd3<=6;bcd2<=7;bcd1<=0;bcd0<=5; end
			6706: begin bcd3<=6;bcd2<=7;bcd1<=0;bcd0<=6; end
			6707: begin bcd3<=6;bcd2<=7;bcd1<=0;bcd0<=7; end
			6708: begin bcd3<=6;bcd2<=7;bcd1<=0;bcd0<=8; end
			6709: begin bcd3<=6;bcd2<=7;bcd1<=0;bcd0<=9; end
			6710: begin bcd3<=6;bcd2<=7;bcd1<=1;bcd0<=0; end
			6711: begin bcd3<=6;bcd2<=7;bcd1<=1;bcd0<=1; end
			6712: begin bcd3<=6;bcd2<=7;bcd1<=1;bcd0<=2; end
			6713: begin bcd3<=6;bcd2<=7;bcd1<=1;bcd0<=3; end
			6714: begin bcd3<=6;bcd2<=7;bcd1<=1;bcd0<=4; end
			6715: begin bcd3<=6;bcd2<=7;bcd1<=1;bcd0<=5; end
			6716: begin bcd3<=6;bcd2<=7;bcd1<=1;bcd0<=6; end
			6717: begin bcd3<=6;bcd2<=7;bcd1<=1;bcd0<=7; end
			6718: begin bcd3<=6;bcd2<=7;bcd1<=1;bcd0<=8; end
			6719: begin bcd3<=6;bcd2<=7;bcd1<=1;bcd0<=9; end
			6720: begin bcd3<=6;bcd2<=7;bcd1<=2;bcd0<=0; end
			6721: begin bcd3<=6;bcd2<=7;bcd1<=2;bcd0<=1; end
			6722: begin bcd3<=6;bcd2<=7;bcd1<=2;bcd0<=2; end
			6723: begin bcd3<=6;bcd2<=7;bcd1<=2;bcd0<=3; end
			6724: begin bcd3<=6;bcd2<=7;bcd1<=2;bcd0<=4; end
			6725: begin bcd3<=6;bcd2<=7;bcd1<=2;bcd0<=5; end
			6726: begin bcd3<=6;bcd2<=7;bcd1<=2;bcd0<=6; end
			6727: begin bcd3<=6;bcd2<=7;bcd1<=2;bcd0<=7; end
			6728: begin bcd3<=6;bcd2<=7;bcd1<=2;bcd0<=8; end
			6729: begin bcd3<=6;bcd2<=7;bcd1<=2;bcd0<=9; end
			6730: begin bcd3<=6;bcd2<=7;bcd1<=3;bcd0<=0; end
			6731: begin bcd3<=6;bcd2<=7;bcd1<=3;bcd0<=1; end
			6732: begin bcd3<=6;bcd2<=7;bcd1<=3;bcd0<=2; end
			6733: begin bcd3<=6;bcd2<=7;bcd1<=3;bcd0<=3; end
			6734: begin bcd3<=6;bcd2<=7;bcd1<=3;bcd0<=4; end
			6735: begin bcd3<=6;bcd2<=7;bcd1<=3;bcd0<=5; end
			6736: begin bcd3<=6;bcd2<=7;bcd1<=3;bcd0<=6; end
			6737: begin bcd3<=6;bcd2<=7;bcd1<=3;bcd0<=7; end
			6738: begin bcd3<=6;bcd2<=7;bcd1<=3;bcd0<=8; end
			6739: begin bcd3<=6;bcd2<=7;bcd1<=3;bcd0<=9; end
			6740: begin bcd3<=6;bcd2<=7;bcd1<=4;bcd0<=0; end
			6741: begin bcd3<=6;bcd2<=7;bcd1<=4;bcd0<=1; end
			6742: begin bcd3<=6;bcd2<=7;bcd1<=4;bcd0<=2; end
			6743: begin bcd3<=6;bcd2<=7;bcd1<=4;bcd0<=3; end
			6744: begin bcd3<=6;bcd2<=7;bcd1<=4;bcd0<=4; end
			6745: begin bcd3<=6;bcd2<=7;bcd1<=4;bcd0<=5; end
			6746: begin bcd3<=6;bcd2<=7;bcd1<=4;bcd0<=6; end
			6747: begin bcd3<=6;bcd2<=7;bcd1<=4;bcd0<=7; end
			6748: begin bcd3<=6;bcd2<=7;bcd1<=4;bcd0<=8; end
			6749: begin bcd3<=6;bcd2<=7;bcd1<=4;bcd0<=9; end
			6750: begin bcd3<=6;bcd2<=7;bcd1<=5;bcd0<=0; end
			6751: begin bcd3<=6;bcd2<=7;bcd1<=5;bcd0<=1; end
			6752: begin bcd3<=6;bcd2<=7;bcd1<=5;bcd0<=2; end
			6753: begin bcd3<=6;bcd2<=7;bcd1<=5;bcd0<=3; end
			6754: begin bcd3<=6;bcd2<=7;bcd1<=5;bcd0<=4; end
			6755: begin bcd3<=6;bcd2<=7;bcd1<=5;bcd0<=5; end
			6756: begin bcd3<=6;bcd2<=7;bcd1<=5;bcd0<=6; end
			6757: begin bcd3<=6;bcd2<=7;bcd1<=5;bcd0<=7; end
			6758: begin bcd3<=6;bcd2<=7;bcd1<=5;bcd0<=8; end
			6759: begin bcd3<=6;bcd2<=7;bcd1<=5;bcd0<=9; end
			6760: begin bcd3<=6;bcd2<=7;bcd1<=6;bcd0<=0; end
			6761: begin bcd3<=6;bcd2<=7;bcd1<=6;bcd0<=1; end
			6762: begin bcd3<=6;bcd2<=7;bcd1<=6;bcd0<=2; end
			6763: begin bcd3<=6;bcd2<=7;bcd1<=6;bcd0<=3; end
			6764: begin bcd3<=6;bcd2<=7;bcd1<=6;bcd0<=4; end
			6765: begin bcd3<=6;bcd2<=7;bcd1<=6;bcd0<=5; end
			6766: begin bcd3<=6;bcd2<=7;bcd1<=6;bcd0<=6; end
			6767: begin bcd3<=6;bcd2<=7;bcd1<=6;bcd0<=7; end
			6768: begin bcd3<=6;bcd2<=7;bcd1<=6;bcd0<=8; end
			6769: begin bcd3<=6;bcd2<=7;bcd1<=6;bcd0<=9; end
			6770: begin bcd3<=6;bcd2<=7;bcd1<=7;bcd0<=0; end
			6771: begin bcd3<=6;bcd2<=7;bcd1<=7;bcd0<=1; end
			6772: begin bcd3<=6;bcd2<=7;bcd1<=7;bcd0<=2; end
			6773: begin bcd3<=6;bcd2<=7;bcd1<=7;bcd0<=3; end
			6774: begin bcd3<=6;bcd2<=7;bcd1<=7;bcd0<=4; end
			6775: begin bcd3<=6;bcd2<=7;bcd1<=7;bcd0<=5; end
			6776: begin bcd3<=6;bcd2<=7;bcd1<=7;bcd0<=6; end
			6777: begin bcd3<=6;bcd2<=7;bcd1<=7;bcd0<=7; end
			6778: begin bcd3<=6;bcd2<=7;bcd1<=7;bcd0<=8; end
			6779: begin bcd3<=6;bcd2<=7;bcd1<=7;bcd0<=9; end
			6780: begin bcd3<=6;bcd2<=7;bcd1<=8;bcd0<=0; end
			6781: begin bcd3<=6;bcd2<=7;bcd1<=8;bcd0<=1; end
			6782: begin bcd3<=6;bcd2<=7;bcd1<=8;bcd0<=2; end
			6783: begin bcd3<=6;bcd2<=7;bcd1<=8;bcd0<=3; end
			6784: begin bcd3<=6;bcd2<=7;bcd1<=8;bcd0<=4; end
			6785: begin bcd3<=6;bcd2<=7;bcd1<=8;bcd0<=5; end
			6786: begin bcd3<=6;bcd2<=7;bcd1<=8;bcd0<=6; end
			6787: begin bcd3<=6;bcd2<=7;bcd1<=8;bcd0<=7; end
			6788: begin bcd3<=6;bcd2<=7;bcd1<=8;bcd0<=8; end
			6789: begin bcd3<=6;bcd2<=7;bcd1<=8;bcd0<=9; end
			6790: begin bcd3<=6;bcd2<=7;bcd1<=9;bcd0<=0; end
			6791: begin bcd3<=6;bcd2<=7;bcd1<=9;bcd0<=1; end
			6792: begin bcd3<=6;bcd2<=7;bcd1<=9;bcd0<=2; end
			6793: begin bcd3<=6;bcd2<=7;bcd1<=9;bcd0<=3; end
			6794: begin bcd3<=6;bcd2<=7;bcd1<=9;bcd0<=4; end
			6795: begin bcd3<=6;bcd2<=7;bcd1<=9;bcd0<=5; end
			6796: begin bcd3<=6;bcd2<=7;bcd1<=9;bcd0<=6; end
			6797: begin bcd3<=6;bcd2<=7;bcd1<=9;bcd0<=7; end
			6798: begin bcd3<=6;bcd2<=7;bcd1<=9;bcd0<=8; end
			6799: begin bcd3<=6;bcd2<=7;bcd1<=9;bcd0<=9; end
			6800: begin bcd3<=6;bcd2<=8;bcd1<=0;bcd0<=0; end
			6801: begin bcd3<=6;bcd2<=8;bcd1<=0;bcd0<=1; end
			6802: begin bcd3<=6;bcd2<=8;bcd1<=0;bcd0<=2; end
			6803: begin bcd3<=6;bcd2<=8;bcd1<=0;bcd0<=3; end
			6804: begin bcd3<=6;bcd2<=8;bcd1<=0;bcd0<=4; end
			6805: begin bcd3<=6;bcd2<=8;bcd1<=0;bcd0<=5; end
			6806: begin bcd3<=6;bcd2<=8;bcd1<=0;bcd0<=6; end
			6807: begin bcd3<=6;bcd2<=8;bcd1<=0;bcd0<=7; end
			6808: begin bcd3<=6;bcd2<=8;bcd1<=0;bcd0<=8; end
			6809: begin bcd3<=6;bcd2<=8;bcd1<=0;bcd0<=9; end
			6810: begin bcd3<=6;bcd2<=8;bcd1<=1;bcd0<=0; end
			6811: begin bcd3<=6;bcd2<=8;bcd1<=1;bcd0<=1; end
			6812: begin bcd3<=6;bcd2<=8;bcd1<=1;bcd0<=2; end
			6813: begin bcd3<=6;bcd2<=8;bcd1<=1;bcd0<=3; end
			6814: begin bcd3<=6;bcd2<=8;bcd1<=1;bcd0<=4; end
			6815: begin bcd3<=6;bcd2<=8;bcd1<=1;bcd0<=5; end
			6816: begin bcd3<=6;bcd2<=8;bcd1<=1;bcd0<=6; end
			6817: begin bcd3<=6;bcd2<=8;bcd1<=1;bcd0<=7; end
			6818: begin bcd3<=6;bcd2<=8;bcd1<=1;bcd0<=8; end
			6819: begin bcd3<=6;bcd2<=8;bcd1<=1;bcd0<=9; end
			6820: begin bcd3<=6;bcd2<=8;bcd1<=2;bcd0<=0; end
			6821: begin bcd3<=6;bcd2<=8;bcd1<=2;bcd0<=1; end
			6822: begin bcd3<=6;bcd2<=8;bcd1<=2;bcd0<=2; end
			6823: begin bcd3<=6;bcd2<=8;bcd1<=2;bcd0<=3; end
			6824: begin bcd3<=6;bcd2<=8;bcd1<=2;bcd0<=4; end
			6825: begin bcd3<=6;bcd2<=8;bcd1<=2;bcd0<=5; end
			6826: begin bcd3<=6;bcd2<=8;bcd1<=2;bcd0<=6; end
			6827: begin bcd3<=6;bcd2<=8;bcd1<=2;bcd0<=7; end
			6828: begin bcd3<=6;bcd2<=8;bcd1<=2;bcd0<=8; end
			6829: begin bcd3<=6;bcd2<=8;bcd1<=2;bcd0<=9; end
			6830: begin bcd3<=6;bcd2<=8;bcd1<=3;bcd0<=0; end
			6831: begin bcd3<=6;bcd2<=8;bcd1<=3;bcd0<=1; end
			6832: begin bcd3<=6;bcd2<=8;bcd1<=3;bcd0<=2; end
			6833: begin bcd3<=6;bcd2<=8;bcd1<=3;bcd0<=3; end
			6834: begin bcd3<=6;bcd2<=8;bcd1<=3;bcd0<=4; end
			6835: begin bcd3<=6;bcd2<=8;bcd1<=3;bcd0<=5; end
			6836: begin bcd3<=6;bcd2<=8;bcd1<=3;bcd0<=6; end
			6837: begin bcd3<=6;bcd2<=8;bcd1<=3;bcd0<=7; end
			6838: begin bcd3<=6;bcd2<=8;bcd1<=3;bcd0<=8; end
			6839: begin bcd3<=6;bcd2<=8;bcd1<=3;bcd0<=9; end
			6840: begin bcd3<=6;bcd2<=8;bcd1<=4;bcd0<=0; end
			6841: begin bcd3<=6;bcd2<=8;bcd1<=4;bcd0<=1; end
			6842: begin bcd3<=6;bcd2<=8;bcd1<=4;bcd0<=2; end
			6843: begin bcd3<=6;bcd2<=8;bcd1<=4;bcd0<=3; end
			6844: begin bcd3<=6;bcd2<=8;bcd1<=4;bcd0<=4; end
			6845: begin bcd3<=6;bcd2<=8;bcd1<=4;bcd0<=5; end
			6846: begin bcd3<=6;bcd2<=8;bcd1<=4;bcd0<=6; end
			6847: begin bcd3<=6;bcd2<=8;bcd1<=4;bcd0<=7; end
			6848: begin bcd3<=6;bcd2<=8;bcd1<=4;bcd0<=8; end
			6849: begin bcd3<=6;bcd2<=8;bcd1<=4;bcd0<=9; end
			6850: begin bcd3<=6;bcd2<=8;bcd1<=5;bcd0<=0; end
			6851: begin bcd3<=6;bcd2<=8;bcd1<=5;bcd0<=1; end
			6852: begin bcd3<=6;bcd2<=8;bcd1<=5;bcd0<=2; end
			6853: begin bcd3<=6;bcd2<=8;bcd1<=5;bcd0<=3; end
			6854: begin bcd3<=6;bcd2<=8;bcd1<=5;bcd0<=4; end
			6855: begin bcd3<=6;bcd2<=8;bcd1<=5;bcd0<=5; end
			6856: begin bcd3<=6;bcd2<=8;bcd1<=5;bcd0<=6; end
			6857: begin bcd3<=6;bcd2<=8;bcd1<=5;bcd0<=7; end
			6858: begin bcd3<=6;bcd2<=8;bcd1<=5;bcd0<=8; end
			6859: begin bcd3<=6;bcd2<=8;bcd1<=5;bcd0<=9; end
			6860: begin bcd3<=6;bcd2<=8;bcd1<=6;bcd0<=0; end
			6861: begin bcd3<=6;bcd2<=8;bcd1<=6;bcd0<=1; end
			6862: begin bcd3<=6;bcd2<=8;bcd1<=6;bcd0<=2; end
			6863: begin bcd3<=6;bcd2<=8;bcd1<=6;bcd0<=3; end
			6864: begin bcd3<=6;bcd2<=8;bcd1<=6;bcd0<=4; end
			6865: begin bcd3<=6;bcd2<=8;bcd1<=6;bcd0<=5; end
			6866: begin bcd3<=6;bcd2<=8;bcd1<=6;bcd0<=6; end
			6867: begin bcd3<=6;bcd2<=8;bcd1<=6;bcd0<=7; end
			6868: begin bcd3<=6;bcd2<=8;bcd1<=6;bcd0<=8; end
			6869: begin bcd3<=6;bcd2<=8;bcd1<=6;bcd0<=9; end
			6870: begin bcd3<=6;bcd2<=8;bcd1<=7;bcd0<=0; end
			6871: begin bcd3<=6;bcd2<=8;bcd1<=7;bcd0<=1; end
			6872: begin bcd3<=6;bcd2<=8;bcd1<=7;bcd0<=2; end
			6873: begin bcd3<=6;bcd2<=8;bcd1<=7;bcd0<=3; end
			6874: begin bcd3<=6;bcd2<=8;bcd1<=7;bcd0<=4; end
			6875: begin bcd3<=6;bcd2<=8;bcd1<=7;bcd0<=5; end
			6876: begin bcd3<=6;bcd2<=8;bcd1<=7;bcd0<=6; end
			6877: begin bcd3<=6;bcd2<=8;bcd1<=7;bcd0<=7; end
			6878: begin bcd3<=6;bcd2<=8;bcd1<=7;bcd0<=8; end
			6879: begin bcd3<=6;bcd2<=8;bcd1<=7;bcd0<=9; end
			6880: begin bcd3<=6;bcd2<=8;bcd1<=8;bcd0<=0; end
			6881: begin bcd3<=6;bcd2<=8;bcd1<=8;bcd0<=1; end
			6882: begin bcd3<=6;bcd2<=8;bcd1<=8;bcd0<=2; end
			6883: begin bcd3<=6;bcd2<=8;bcd1<=8;bcd0<=3; end
			6884: begin bcd3<=6;bcd2<=8;bcd1<=8;bcd0<=4; end
			6885: begin bcd3<=6;bcd2<=8;bcd1<=8;bcd0<=5; end
			6886: begin bcd3<=6;bcd2<=8;bcd1<=8;bcd0<=6; end
			6887: begin bcd3<=6;bcd2<=8;bcd1<=8;bcd0<=7; end
			6888: begin bcd3<=6;bcd2<=8;bcd1<=8;bcd0<=8; end
			6889: begin bcd3<=6;bcd2<=8;bcd1<=8;bcd0<=9; end
			6890: begin bcd3<=6;bcd2<=8;bcd1<=9;bcd0<=0; end
			6891: begin bcd3<=6;bcd2<=8;bcd1<=9;bcd0<=1; end
			6892: begin bcd3<=6;bcd2<=8;bcd1<=9;bcd0<=2; end
			6893: begin bcd3<=6;bcd2<=8;bcd1<=9;bcd0<=3; end
			6894: begin bcd3<=6;bcd2<=8;bcd1<=9;bcd0<=4; end
			6895: begin bcd3<=6;bcd2<=8;bcd1<=9;bcd0<=5; end
			6896: begin bcd3<=6;bcd2<=8;bcd1<=9;bcd0<=6; end
			6897: begin bcd3<=6;bcd2<=8;bcd1<=9;bcd0<=7; end
			6898: begin bcd3<=6;bcd2<=8;bcd1<=9;bcd0<=8; end
			6899: begin bcd3<=6;bcd2<=8;bcd1<=9;bcd0<=9; end
			6900: begin bcd3<=6;bcd2<=9;bcd1<=0;bcd0<=0; end
			6901: begin bcd3<=6;bcd2<=9;bcd1<=0;bcd0<=1; end
			6902: begin bcd3<=6;bcd2<=9;bcd1<=0;bcd0<=2; end
			6903: begin bcd3<=6;bcd2<=9;bcd1<=0;bcd0<=3; end
			6904: begin bcd3<=6;bcd2<=9;bcd1<=0;bcd0<=4; end
			6905: begin bcd3<=6;bcd2<=9;bcd1<=0;bcd0<=5; end
			6906: begin bcd3<=6;bcd2<=9;bcd1<=0;bcd0<=6; end
			6907: begin bcd3<=6;bcd2<=9;bcd1<=0;bcd0<=7; end
			6908: begin bcd3<=6;bcd2<=9;bcd1<=0;bcd0<=8; end
			6909: begin bcd3<=6;bcd2<=9;bcd1<=0;bcd0<=9; end
			6910: begin bcd3<=6;bcd2<=9;bcd1<=1;bcd0<=0; end
			6911: begin bcd3<=6;bcd2<=9;bcd1<=1;bcd0<=1; end
			6912: begin bcd3<=6;bcd2<=9;bcd1<=1;bcd0<=2; end
			6913: begin bcd3<=6;bcd2<=9;bcd1<=1;bcd0<=3; end
			6914: begin bcd3<=6;bcd2<=9;bcd1<=1;bcd0<=4; end
			6915: begin bcd3<=6;bcd2<=9;bcd1<=1;bcd0<=5; end
			6916: begin bcd3<=6;bcd2<=9;bcd1<=1;bcd0<=6; end
			6917: begin bcd3<=6;bcd2<=9;bcd1<=1;bcd0<=7; end
			6918: begin bcd3<=6;bcd2<=9;bcd1<=1;bcd0<=8; end
			6919: begin bcd3<=6;bcd2<=9;bcd1<=1;bcd0<=9; end
			6920: begin bcd3<=6;bcd2<=9;bcd1<=2;bcd0<=0; end
			6921: begin bcd3<=6;bcd2<=9;bcd1<=2;bcd0<=1; end
			6922: begin bcd3<=6;bcd2<=9;bcd1<=2;bcd0<=2; end
			6923: begin bcd3<=6;bcd2<=9;bcd1<=2;bcd0<=3; end
			6924: begin bcd3<=6;bcd2<=9;bcd1<=2;bcd0<=4; end
			6925: begin bcd3<=6;bcd2<=9;bcd1<=2;bcd0<=5; end
			6926: begin bcd3<=6;bcd2<=9;bcd1<=2;bcd0<=6; end
			6927: begin bcd3<=6;bcd2<=9;bcd1<=2;bcd0<=7; end
			6928: begin bcd3<=6;bcd2<=9;bcd1<=2;bcd0<=8; end
			6929: begin bcd3<=6;bcd2<=9;bcd1<=2;bcd0<=9; end
			6930: begin bcd3<=6;bcd2<=9;bcd1<=3;bcd0<=0; end
			6931: begin bcd3<=6;bcd2<=9;bcd1<=3;bcd0<=1; end
			6932: begin bcd3<=6;bcd2<=9;bcd1<=3;bcd0<=2; end
			6933: begin bcd3<=6;bcd2<=9;bcd1<=3;bcd0<=3; end
			6934: begin bcd3<=6;bcd2<=9;bcd1<=3;bcd0<=4; end
			6935: begin bcd3<=6;bcd2<=9;bcd1<=3;bcd0<=5; end
			6936: begin bcd3<=6;bcd2<=9;bcd1<=3;bcd0<=6; end
			6937: begin bcd3<=6;bcd2<=9;bcd1<=3;bcd0<=7; end
			6938: begin bcd3<=6;bcd2<=9;bcd1<=3;bcd0<=8; end
			6939: begin bcd3<=6;bcd2<=9;bcd1<=3;bcd0<=9; end
			6940: begin bcd3<=6;bcd2<=9;bcd1<=4;bcd0<=0; end
			6941: begin bcd3<=6;bcd2<=9;bcd1<=4;bcd0<=1; end
			6942: begin bcd3<=6;bcd2<=9;bcd1<=4;bcd0<=2; end
			6943: begin bcd3<=6;bcd2<=9;bcd1<=4;bcd0<=3; end
			6944: begin bcd3<=6;bcd2<=9;bcd1<=4;bcd0<=4; end
			6945: begin bcd3<=6;bcd2<=9;bcd1<=4;bcd0<=5; end
			6946: begin bcd3<=6;bcd2<=9;bcd1<=4;bcd0<=6; end
			6947: begin bcd3<=6;bcd2<=9;bcd1<=4;bcd0<=7; end
			6948: begin bcd3<=6;bcd2<=9;bcd1<=4;bcd0<=8; end
			6949: begin bcd3<=6;bcd2<=9;bcd1<=4;bcd0<=9; end
			6950: begin bcd3<=6;bcd2<=9;bcd1<=5;bcd0<=0; end
			6951: begin bcd3<=6;bcd2<=9;bcd1<=5;bcd0<=1; end
			6952: begin bcd3<=6;bcd2<=9;bcd1<=5;bcd0<=2; end
			6953: begin bcd3<=6;bcd2<=9;bcd1<=5;bcd0<=3; end
			6954: begin bcd3<=6;bcd2<=9;bcd1<=5;bcd0<=4; end
			6955: begin bcd3<=6;bcd2<=9;bcd1<=5;bcd0<=5; end
			6956: begin bcd3<=6;bcd2<=9;bcd1<=5;bcd0<=6; end
			6957: begin bcd3<=6;bcd2<=9;bcd1<=5;bcd0<=7; end
			6958: begin bcd3<=6;bcd2<=9;bcd1<=5;bcd0<=8; end
			6959: begin bcd3<=6;bcd2<=9;bcd1<=5;bcd0<=9; end
			6960: begin bcd3<=6;bcd2<=9;bcd1<=6;bcd0<=0; end
			6961: begin bcd3<=6;bcd2<=9;bcd1<=6;bcd0<=1; end
			6962: begin bcd3<=6;bcd2<=9;bcd1<=6;bcd0<=2; end
			6963: begin bcd3<=6;bcd2<=9;bcd1<=6;bcd0<=3; end
			6964: begin bcd3<=6;bcd2<=9;bcd1<=6;bcd0<=4; end
			6965: begin bcd3<=6;bcd2<=9;bcd1<=6;bcd0<=5; end
			6966: begin bcd3<=6;bcd2<=9;bcd1<=6;bcd0<=6; end
			6967: begin bcd3<=6;bcd2<=9;bcd1<=6;bcd0<=7; end
			6968: begin bcd3<=6;bcd2<=9;bcd1<=6;bcd0<=8; end
			6969: begin bcd3<=6;bcd2<=9;bcd1<=6;bcd0<=9; end
			6970: begin bcd3<=6;bcd2<=9;bcd1<=7;bcd0<=0; end
			6971: begin bcd3<=6;bcd2<=9;bcd1<=7;bcd0<=1; end
			6972: begin bcd3<=6;bcd2<=9;bcd1<=7;bcd0<=2; end
			6973: begin bcd3<=6;bcd2<=9;bcd1<=7;bcd0<=3; end
			6974: begin bcd3<=6;bcd2<=9;bcd1<=7;bcd0<=4; end
			6975: begin bcd3<=6;bcd2<=9;bcd1<=7;bcd0<=5; end
			6976: begin bcd3<=6;bcd2<=9;bcd1<=7;bcd0<=6; end
			6977: begin bcd3<=6;bcd2<=9;bcd1<=7;bcd0<=7; end
			6978: begin bcd3<=6;bcd2<=9;bcd1<=7;bcd0<=8; end
			6979: begin bcd3<=6;bcd2<=9;bcd1<=7;bcd0<=9; end
			6980: begin bcd3<=6;bcd2<=9;bcd1<=8;bcd0<=0; end
			6981: begin bcd3<=6;bcd2<=9;bcd1<=8;bcd0<=1; end
			6982: begin bcd3<=6;bcd2<=9;bcd1<=8;bcd0<=2; end
			6983: begin bcd3<=6;bcd2<=9;bcd1<=8;bcd0<=3; end
			6984: begin bcd3<=6;bcd2<=9;bcd1<=8;bcd0<=4; end
			6985: begin bcd3<=6;bcd2<=9;bcd1<=8;bcd0<=5; end
			6986: begin bcd3<=6;bcd2<=9;bcd1<=8;bcd0<=6; end
			6987: begin bcd3<=6;bcd2<=9;bcd1<=8;bcd0<=7; end
			6988: begin bcd3<=6;bcd2<=9;bcd1<=8;bcd0<=8; end
			6989: begin bcd3<=6;bcd2<=9;bcd1<=8;bcd0<=9; end
			6990: begin bcd3<=6;bcd2<=9;bcd1<=9;bcd0<=0; end
			6991: begin bcd3<=6;bcd2<=9;bcd1<=9;bcd0<=1; end
			6992: begin bcd3<=6;bcd2<=9;bcd1<=9;bcd0<=2; end
			6993: begin bcd3<=6;bcd2<=9;bcd1<=9;bcd0<=3; end
			6994: begin bcd3<=6;bcd2<=9;bcd1<=9;bcd0<=4; end
			6995: begin bcd3<=6;bcd2<=9;bcd1<=9;bcd0<=5; end
			6996: begin bcd3<=6;bcd2<=9;bcd1<=9;bcd0<=6; end
			6997: begin bcd3<=6;bcd2<=9;bcd1<=9;bcd0<=7; end
			6998: begin bcd3<=6;bcd2<=9;bcd1<=9;bcd0<=8; end
			6999: begin bcd3<=6;bcd2<=9;bcd1<=9;bcd0<=9; end
			7000: begin bcd3<=7;bcd2<=0;bcd1<=0;bcd0<=0; end
			7001: begin bcd3<=7;bcd2<=0;bcd1<=0;bcd0<=1; end
			7002: begin bcd3<=7;bcd2<=0;bcd1<=0;bcd0<=2; end
			7003: begin bcd3<=7;bcd2<=0;bcd1<=0;bcd0<=3; end
			7004: begin bcd3<=7;bcd2<=0;bcd1<=0;bcd0<=4; end
			7005: begin bcd3<=7;bcd2<=0;bcd1<=0;bcd0<=5; end
			7006: begin bcd3<=7;bcd2<=0;bcd1<=0;bcd0<=6; end
			7007: begin bcd3<=7;bcd2<=0;bcd1<=0;bcd0<=7; end
			7008: begin bcd3<=7;bcd2<=0;bcd1<=0;bcd0<=8; end
			7009: begin bcd3<=7;bcd2<=0;bcd1<=0;bcd0<=9; end
			7010: begin bcd3<=7;bcd2<=0;bcd1<=1;bcd0<=0; end
			7011: begin bcd3<=7;bcd2<=0;bcd1<=1;bcd0<=1; end
			7012: begin bcd3<=7;bcd2<=0;bcd1<=1;bcd0<=2; end
			7013: begin bcd3<=7;bcd2<=0;bcd1<=1;bcd0<=3; end
			7014: begin bcd3<=7;bcd2<=0;bcd1<=1;bcd0<=4; end
			7015: begin bcd3<=7;bcd2<=0;bcd1<=1;bcd0<=5; end
			7016: begin bcd3<=7;bcd2<=0;bcd1<=1;bcd0<=6; end
			7017: begin bcd3<=7;bcd2<=0;bcd1<=1;bcd0<=7; end
			7018: begin bcd3<=7;bcd2<=0;bcd1<=1;bcd0<=8; end
			7019: begin bcd3<=7;bcd2<=0;bcd1<=1;bcd0<=9; end
			7020: begin bcd3<=7;bcd2<=0;bcd1<=2;bcd0<=0; end
			7021: begin bcd3<=7;bcd2<=0;bcd1<=2;bcd0<=1; end
			7022: begin bcd3<=7;bcd2<=0;bcd1<=2;bcd0<=2; end
			7023: begin bcd3<=7;bcd2<=0;bcd1<=2;bcd0<=3; end
			7024: begin bcd3<=7;bcd2<=0;bcd1<=2;bcd0<=4; end
			7025: begin bcd3<=7;bcd2<=0;bcd1<=2;bcd0<=5; end
			7026: begin bcd3<=7;bcd2<=0;bcd1<=2;bcd0<=6; end
			7027: begin bcd3<=7;bcd2<=0;bcd1<=2;bcd0<=7; end
			7028: begin bcd3<=7;bcd2<=0;bcd1<=2;bcd0<=8; end
			7029: begin bcd3<=7;bcd2<=0;bcd1<=2;bcd0<=9; end
			7030: begin bcd3<=7;bcd2<=0;bcd1<=3;bcd0<=0; end
			7031: begin bcd3<=7;bcd2<=0;bcd1<=3;bcd0<=1; end
			7032: begin bcd3<=7;bcd2<=0;bcd1<=3;bcd0<=2; end
			7033: begin bcd3<=7;bcd2<=0;bcd1<=3;bcd0<=3; end
			7034: begin bcd3<=7;bcd2<=0;bcd1<=3;bcd0<=4; end
			7035: begin bcd3<=7;bcd2<=0;bcd1<=3;bcd0<=5; end
			7036: begin bcd3<=7;bcd2<=0;bcd1<=3;bcd0<=6; end
			7037: begin bcd3<=7;bcd2<=0;bcd1<=3;bcd0<=7; end
			7038: begin bcd3<=7;bcd2<=0;bcd1<=3;bcd0<=8; end
			7039: begin bcd3<=7;bcd2<=0;bcd1<=3;bcd0<=9; end
			7040: begin bcd3<=7;bcd2<=0;bcd1<=4;bcd0<=0; end
			7041: begin bcd3<=7;bcd2<=0;bcd1<=4;bcd0<=1; end
			7042: begin bcd3<=7;bcd2<=0;bcd1<=4;bcd0<=2; end
			7043: begin bcd3<=7;bcd2<=0;bcd1<=4;bcd0<=3; end
			7044: begin bcd3<=7;bcd2<=0;bcd1<=4;bcd0<=4; end
			7045: begin bcd3<=7;bcd2<=0;bcd1<=4;bcd0<=5; end
			7046: begin bcd3<=7;bcd2<=0;bcd1<=4;bcd0<=6; end
			7047: begin bcd3<=7;bcd2<=0;bcd1<=4;bcd0<=7; end
			7048: begin bcd3<=7;bcd2<=0;bcd1<=4;bcd0<=8; end
			7049: begin bcd3<=7;bcd2<=0;bcd1<=4;bcd0<=9; end
			7050: begin bcd3<=7;bcd2<=0;bcd1<=5;bcd0<=0; end
			7051: begin bcd3<=7;bcd2<=0;bcd1<=5;bcd0<=1; end
			7052: begin bcd3<=7;bcd2<=0;bcd1<=5;bcd0<=2; end
			7053: begin bcd3<=7;bcd2<=0;bcd1<=5;bcd0<=3; end
			7054: begin bcd3<=7;bcd2<=0;bcd1<=5;bcd0<=4; end
			7055: begin bcd3<=7;bcd2<=0;bcd1<=5;bcd0<=5; end
			7056: begin bcd3<=7;bcd2<=0;bcd1<=5;bcd0<=6; end
			7057: begin bcd3<=7;bcd2<=0;bcd1<=5;bcd0<=7; end
			7058: begin bcd3<=7;bcd2<=0;bcd1<=5;bcd0<=8; end
			7059: begin bcd3<=7;bcd2<=0;bcd1<=5;bcd0<=9; end
			7060: begin bcd3<=7;bcd2<=0;bcd1<=6;bcd0<=0; end
			7061: begin bcd3<=7;bcd2<=0;bcd1<=6;bcd0<=1; end
			7062: begin bcd3<=7;bcd2<=0;bcd1<=6;bcd0<=2; end
			7063: begin bcd3<=7;bcd2<=0;bcd1<=6;bcd0<=3; end
			7064: begin bcd3<=7;bcd2<=0;bcd1<=6;bcd0<=4; end
			7065: begin bcd3<=7;bcd2<=0;bcd1<=6;bcd0<=5; end
			7066: begin bcd3<=7;bcd2<=0;bcd1<=6;bcd0<=6; end
			7067: begin bcd3<=7;bcd2<=0;bcd1<=6;bcd0<=7; end
			7068: begin bcd3<=7;bcd2<=0;bcd1<=6;bcd0<=8; end
			7069: begin bcd3<=7;bcd2<=0;bcd1<=6;bcd0<=9; end
			7070: begin bcd3<=7;bcd2<=0;bcd1<=7;bcd0<=0; end
			7071: begin bcd3<=7;bcd2<=0;bcd1<=7;bcd0<=1; end
			7072: begin bcd3<=7;bcd2<=0;bcd1<=7;bcd0<=2; end
			7073: begin bcd3<=7;bcd2<=0;bcd1<=7;bcd0<=3; end
			7074: begin bcd3<=7;bcd2<=0;bcd1<=7;bcd0<=4; end
			7075: begin bcd3<=7;bcd2<=0;bcd1<=7;bcd0<=5; end
			7076: begin bcd3<=7;bcd2<=0;bcd1<=7;bcd0<=6; end
			7077: begin bcd3<=7;bcd2<=0;bcd1<=7;bcd0<=7; end
			7078: begin bcd3<=7;bcd2<=0;bcd1<=7;bcd0<=8; end
			7079: begin bcd3<=7;bcd2<=0;bcd1<=7;bcd0<=9; end
			7080: begin bcd3<=7;bcd2<=0;bcd1<=8;bcd0<=0; end
			7081: begin bcd3<=7;bcd2<=0;bcd1<=8;bcd0<=1; end
			7082: begin bcd3<=7;bcd2<=0;bcd1<=8;bcd0<=2; end
			7083: begin bcd3<=7;bcd2<=0;bcd1<=8;bcd0<=3; end
			7084: begin bcd3<=7;bcd2<=0;bcd1<=8;bcd0<=4; end
			7085: begin bcd3<=7;bcd2<=0;bcd1<=8;bcd0<=5; end
			7086: begin bcd3<=7;bcd2<=0;bcd1<=8;bcd0<=6; end
			7087: begin bcd3<=7;bcd2<=0;bcd1<=8;bcd0<=7; end
			7088: begin bcd3<=7;bcd2<=0;bcd1<=8;bcd0<=8; end
			7089: begin bcd3<=7;bcd2<=0;bcd1<=8;bcd0<=9; end
			7090: begin bcd3<=7;bcd2<=0;bcd1<=9;bcd0<=0; end
			7091: begin bcd3<=7;bcd2<=0;bcd1<=9;bcd0<=1; end
			7092: begin bcd3<=7;bcd2<=0;bcd1<=9;bcd0<=2; end
			7093: begin bcd3<=7;bcd2<=0;bcd1<=9;bcd0<=3; end
			7094: begin bcd3<=7;bcd2<=0;bcd1<=9;bcd0<=4; end
			7095: begin bcd3<=7;bcd2<=0;bcd1<=9;bcd0<=5; end
			7096: begin bcd3<=7;bcd2<=0;bcd1<=9;bcd0<=6; end
			7097: begin bcd3<=7;bcd2<=0;bcd1<=9;bcd0<=7; end
			7098: begin bcd3<=7;bcd2<=0;bcd1<=9;bcd0<=8; end
			7099: begin bcd3<=7;bcd2<=0;bcd1<=9;bcd0<=9; end
			7100: begin bcd3<=7;bcd2<=1;bcd1<=0;bcd0<=0; end
			7101: begin bcd3<=7;bcd2<=1;bcd1<=0;bcd0<=1; end
			7102: begin bcd3<=7;bcd2<=1;bcd1<=0;bcd0<=2; end
			7103: begin bcd3<=7;bcd2<=1;bcd1<=0;bcd0<=3; end
			7104: begin bcd3<=7;bcd2<=1;bcd1<=0;bcd0<=4; end
			7105: begin bcd3<=7;bcd2<=1;bcd1<=0;bcd0<=5; end
			7106: begin bcd3<=7;bcd2<=1;bcd1<=0;bcd0<=6; end
			7107: begin bcd3<=7;bcd2<=1;bcd1<=0;bcd0<=7; end
			7108: begin bcd3<=7;bcd2<=1;bcd1<=0;bcd0<=8; end
			7109: begin bcd3<=7;bcd2<=1;bcd1<=0;bcd0<=9; end
			7110: begin bcd3<=7;bcd2<=1;bcd1<=1;bcd0<=0; end
			7111: begin bcd3<=7;bcd2<=1;bcd1<=1;bcd0<=1; end
			7112: begin bcd3<=7;bcd2<=1;bcd1<=1;bcd0<=2; end
			7113: begin bcd3<=7;bcd2<=1;bcd1<=1;bcd0<=3; end
			7114: begin bcd3<=7;bcd2<=1;bcd1<=1;bcd0<=4; end
			7115: begin bcd3<=7;bcd2<=1;bcd1<=1;bcd0<=5; end
			7116: begin bcd3<=7;bcd2<=1;bcd1<=1;bcd0<=6; end
			7117: begin bcd3<=7;bcd2<=1;bcd1<=1;bcd0<=7; end
			7118: begin bcd3<=7;bcd2<=1;bcd1<=1;bcd0<=8; end
			7119: begin bcd3<=7;bcd2<=1;bcd1<=1;bcd0<=9; end
			7120: begin bcd3<=7;bcd2<=1;bcd1<=2;bcd0<=0; end
			7121: begin bcd3<=7;bcd2<=1;bcd1<=2;bcd0<=1; end
			7122: begin bcd3<=7;bcd2<=1;bcd1<=2;bcd0<=2; end
			7123: begin bcd3<=7;bcd2<=1;bcd1<=2;bcd0<=3; end
			7124: begin bcd3<=7;bcd2<=1;bcd1<=2;bcd0<=4; end
			7125: begin bcd3<=7;bcd2<=1;bcd1<=2;bcd0<=5; end
			7126: begin bcd3<=7;bcd2<=1;bcd1<=2;bcd0<=6; end
			7127: begin bcd3<=7;bcd2<=1;bcd1<=2;bcd0<=7; end
			7128: begin bcd3<=7;bcd2<=1;bcd1<=2;bcd0<=8; end
			7129: begin bcd3<=7;bcd2<=1;bcd1<=2;bcd0<=9; end
			7130: begin bcd3<=7;bcd2<=1;bcd1<=3;bcd0<=0; end
			7131: begin bcd3<=7;bcd2<=1;bcd1<=3;bcd0<=1; end
			7132: begin bcd3<=7;bcd2<=1;bcd1<=3;bcd0<=2; end
			7133: begin bcd3<=7;bcd2<=1;bcd1<=3;bcd0<=3; end
			7134: begin bcd3<=7;bcd2<=1;bcd1<=3;bcd0<=4; end
			7135: begin bcd3<=7;bcd2<=1;bcd1<=3;bcd0<=5; end
			7136: begin bcd3<=7;bcd2<=1;bcd1<=3;bcd0<=6; end
			7137: begin bcd3<=7;bcd2<=1;bcd1<=3;bcd0<=7; end
			7138: begin bcd3<=7;bcd2<=1;bcd1<=3;bcd0<=8; end
			7139: begin bcd3<=7;bcd2<=1;bcd1<=3;bcd0<=9; end
			7140: begin bcd3<=7;bcd2<=1;bcd1<=4;bcd0<=0; end
			7141: begin bcd3<=7;bcd2<=1;bcd1<=4;bcd0<=1; end
			7142: begin bcd3<=7;bcd2<=1;bcd1<=4;bcd0<=2; end
			7143: begin bcd3<=7;bcd2<=1;bcd1<=4;bcd0<=3; end
			7144: begin bcd3<=7;bcd2<=1;bcd1<=4;bcd0<=4; end
			7145: begin bcd3<=7;bcd2<=1;bcd1<=4;bcd0<=5; end
			7146: begin bcd3<=7;bcd2<=1;bcd1<=4;bcd0<=6; end
			7147: begin bcd3<=7;bcd2<=1;bcd1<=4;bcd0<=7; end
			7148: begin bcd3<=7;bcd2<=1;bcd1<=4;bcd0<=8; end
			7149: begin bcd3<=7;bcd2<=1;bcd1<=4;bcd0<=9; end
			7150: begin bcd3<=7;bcd2<=1;bcd1<=5;bcd0<=0; end
			7151: begin bcd3<=7;bcd2<=1;bcd1<=5;bcd0<=1; end
			7152: begin bcd3<=7;bcd2<=1;bcd1<=5;bcd0<=2; end
			7153: begin bcd3<=7;bcd2<=1;bcd1<=5;bcd0<=3; end
			7154: begin bcd3<=7;bcd2<=1;bcd1<=5;bcd0<=4; end
			7155: begin bcd3<=7;bcd2<=1;bcd1<=5;bcd0<=5; end
			7156: begin bcd3<=7;bcd2<=1;bcd1<=5;bcd0<=6; end
			7157: begin bcd3<=7;bcd2<=1;bcd1<=5;bcd0<=7; end
			7158: begin bcd3<=7;bcd2<=1;bcd1<=5;bcd0<=8; end
			7159: begin bcd3<=7;bcd2<=1;bcd1<=5;bcd0<=9; end
			7160: begin bcd3<=7;bcd2<=1;bcd1<=6;bcd0<=0; end
			7161: begin bcd3<=7;bcd2<=1;bcd1<=6;bcd0<=1; end
			7162: begin bcd3<=7;bcd2<=1;bcd1<=6;bcd0<=2; end
			7163: begin bcd3<=7;bcd2<=1;bcd1<=6;bcd0<=3; end
			7164: begin bcd3<=7;bcd2<=1;bcd1<=6;bcd0<=4; end
			7165: begin bcd3<=7;bcd2<=1;bcd1<=6;bcd0<=5; end
			7166: begin bcd3<=7;bcd2<=1;bcd1<=6;bcd0<=6; end
			7167: begin bcd3<=7;bcd2<=1;bcd1<=6;bcd0<=7; end
			7168: begin bcd3<=7;bcd2<=1;bcd1<=6;bcd0<=8; end
			7169: begin bcd3<=7;bcd2<=1;bcd1<=6;bcd0<=9; end
			7170: begin bcd3<=7;bcd2<=1;bcd1<=7;bcd0<=0; end
			7171: begin bcd3<=7;bcd2<=1;bcd1<=7;bcd0<=1; end
			7172: begin bcd3<=7;bcd2<=1;bcd1<=7;bcd0<=2; end
			7173: begin bcd3<=7;bcd2<=1;bcd1<=7;bcd0<=3; end
			7174: begin bcd3<=7;bcd2<=1;bcd1<=7;bcd0<=4; end
			7175: begin bcd3<=7;bcd2<=1;bcd1<=7;bcd0<=5; end
			7176: begin bcd3<=7;bcd2<=1;bcd1<=7;bcd0<=6; end
			7177: begin bcd3<=7;bcd2<=1;bcd1<=7;bcd0<=7; end
			7178: begin bcd3<=7;bcd2<=1;bcd1<=7;bcd0<=8; end
			7179: begin bcd3<=7;bcd2<=1;bcd1<=7;bcd0<=9; end
			7180: begin bcd3<=7;bcd2<=1;bcd1<=8;bcd0<=0; end
			7181: begin bcd3<=7;bcd2<=1;bcd1<=8;bcd0<=1; end
			7182: begin bcd3<=7;bcd2<=1;bcd1<=8;bcd0<=2; end
			7183: begin bcd3<=7;bcd2<=1;bcd1<=8;bcd0<=3; end
			7184: begin bcd3<=7;bcd2<=1;bcd1<=8;bcd0<=4; end
			7185: begin bcd3<=7;bcd2<=1;bcd1<=8;bcd0<=5; end
			7186: begin bcd3<=7;bcd2<=1;bcd1<=8;bcd0<=6; end
			7187: begin bcd3<=7;bcd2<=1;bcd1<=8;bcd0<=7; end
			7188: begin bcd3<=7;bcd2<=1;bcd1<=8;bcd0<=8; end
			7189: begin bcd3<=7;bcd2<=1;bcd1<=8;bcd0<=9; end
			7190: begin bcd3<=7;bcd2<=1;bcd1<=9;bcd0<=0; end
			7191: begin bcd3<=7;bcd2<=1;bcd1<=9;bcd0<=1; end
			7192: begin bcd3<=7;bcd2<=1;bcd1<=9;bcd0<=2; end
			7193: begin bcd3<=7;bcd2<=1;bcd1<=9;bcd0<=3; end
			7194: begin bcd3<=7;bcd2<=1;bcd1<=9;bcd0<=4; end
			7195: begin bcd3<=7;bcd2<=1;bcd1<=9;bcd0<=5; end
			7196: begin bcd3<=7;bcd2<=1;bcd1<=9;bcd0<=6; end
			7197: begin bcd3<=7;bcd2<=1;bcd1<=9;bcd0<=7; end
			7198: begin bcd3<=7;bcd2<=1;bcd1<=9;bcd0<=8; end
			7199: begin bcd3<=7;bcd2<=1;bcd1<=9;bcd0<=9; end
			7200: begin bcd3<=7;bcd2<=2;bcd1<=0;bcd0<=0; end
			7201: begin bcd3<=7;bcd2<=2;bcd1<=0;bcd0<=1; end
			7202: begin bcd3<=7;bcd2<=2;bcd1<=0;bcd0<=2; end
			7203: begin bcd3<=7;bcd2<=2;bcd1<=0;bcd0<=3; end
			7204: begin bcd3<=7;bcd2<=2;bcd1<=0;bcd0<=4; end
			7205: begin bcd3<=7;bcd2<=2;bcd1<=0;bcd0<=5; end
			7206: begin bcd3<=7;bcd2<=2;bcd1<=0;bcd0<=6; end
			7207: begin bcd3<=7;bcd2<=2;bcd1<=0;bcd0<=7; end
			7208: begin bcd3<=7;bcd2<=2;bcd1<=0;bcd0<=8; end
			7209: begin bcd3<=7;bcd2<=2;bcd1<=0;bcd0<=9; end
			7210: begin bcd3<=7;bcd2<=2;bcd1<=1;bcd0<=0; end
			7211: begin bcd3<=7;bcd2<=2;bcd1<=1;bcd0<=1; end
			7212: begin bcd3<=7;bcd2<=2;bcd1<=1;bcd0<=2; end
			7213: begin bcd3<=7;bcd2<=2;bcd1<=1;bcd0<=3; end
			7214: begin bcd3<=7;bcd2<=2;bcd1<=1;bcd0<=4; end
			7215: begin bcd3<=7;bcd2<=2;bcd1<=1;bcd0<=5; end
			7216: begin bcd3<=7;bcd2<=2;bcd1<=1;bcd0<=6; end
			7217: begin bcd3<=7;bcd2<=2;bcd1<=1;bcd0<=7; end
			7218: begin bcd3<=7;bcd2<=2;bcd1<=1;bcd0<=8; end
			7219: begin bcd3<=7;bcd2<=2;bcd1<=1;bcd0<=9; end
			7220: begin bcd3<=7;bcd2<=2;bcd1<=2;bcd0<=0; end
			7221: begin bcd3<=7;bcd2<=2;bcd1<=2;bcd0<=1; end
			7222: begin bcd3<=7;bcd2<=2;bcd1<=2;bcd0<=2; end
			7223: begin bcd3<=7;bcd2<=2;bcd1<=2;bcd0<=3; end
			7224: begin bcd3<=7;bcd2<=2;bcd1<=2;bcd0<=4; end
			7225: begin bcd3<=7;bcd2<=2;bcd1<=2;bcd0<=5; end
			7226: begin bcd3<=7;bcd2<=2;bcd1<=2;bcd0<=6; end
			7227: begin bcd3<=7;bcd2<=2;bcd1<=2;bcd0<=7; end
			7228: begin bcd3<=7;bcd2<=2;bcd1<=2;bcd0<=8; end
			7229: begin bcd3<=7;bcd2<=2;bcd1<=2;bcd0<=9; end
			7230: begin bcd3<=7;bcd2<=2;bcd1<=3;bcd0<=0; end
			7231: begin bcd3<=7;bcd2<=2;bcd1<=3;bcd0<=1; end
			7232: begin bcd3<=7;bcd2<=2;bcd1<=3;bcd0<=2; end
			7233: begin bcd3<=7;bcd2<=2;bcd1<=3;bcd0<=3; end
			7234: begin bcd3<=7;bcd2<=2;bcd1<=3;bcd0<=4; end
			7235: begin bcd3<=7;bcd2<=2;bcd1<=3;bcd0<=5; end
			7236: begin bcd3<=7;bcd2<=2;bcd1<=3;bcd0<=6; end
			7237: begin bcd3<=7;bcd2<=2;bcd1<=3;bcd0<=7; end
			7238: begin bcd3<=7;bcd2<=2;bcd1<=3;bcd0<=8; end
			7239: begin bcd3<=7;bcd2<=2;bcd1<=3;bcd0<=9; end
			7240: begin bcd3<=7;bcd2<=2;bcd1<=4;bcd0<=0; end
			7241: begin bcd3<=7;bcd2<=2;bcd1<=4;bcd0<=1; end
			7242: begin bcd3<=7;bcd2<=2;bcd1<=4;bcd0<=2; end
			7243: begin bcd3<=7;bcd2<=2;bcd1<=4;bcd0<=3; end
			7244: begin bcd3<=7;bcd2<=2;bcd1<=4;bcd0<=4; end
			7245: begin bcd3<=7;bcd2<=2;bcd1<=4;bcd0<=5; end
			7246: begin bcd3<=7;bcd2<=2;bcd1<=4;bcd0<=6; end
			7247: begin bcd3<=7;bcd2<=2;bcd1<=4;bcd0<=7; end
			7248: begin bcd3<=7;bcd2<=2;bcd1<=4;bcd0<=8; end
			7249: begin bcd3<=7;bcd2<=2;bcd1<=4;bcd0<=9; end
			7250: begin bcd3<=7;bcd2<=2;bcd1<=5;bcd0<=0; end
			7251: begin bcd3<=7;bcd2<=2;bcd1<=5;bcd0<=1; end
			7252: begin bcd3<=7;bcd2<=2;bcd1<=5;bcd0<=2; end
			7253: begin bcd3<=7;bcd2<=2;bcd1<=5;bcd0<=3; end
			7254: begin bcd3<=7;bcd2<=2;bcd1<=5;bcd0<=4; end
			7255: begin bcd3<=7;bcd2<=2;bcd1<=5;bcd0<=5; end
			7256: begin bcd3<=7;bcd2<=2;bcd1<=5;bcd0<=6; end
			7257: begin bcd3<=7;bcd2<=2;bcd1<=5;bcd0<=7; end
			7258: begin bcd3<=7;bcd2<=2;bcd1<=5;bcd0<=8; end
			7259: begin bcd3<=7;bcd2<=2;bcd1<=5;bcd0<=9; end
			7260: begin bcd3<=7;bcd2<=2;bcd1<=6;bcd0<=0; end
			7261: begin bcd3<=7;bcd2<=2;bcd1<=6;bcd0<=1; end
			7262: begin bcd3<=7;bcd2<=2;bcd1<=6;bcd0<=2; end
			7263: begin bcd3<=7;bcd2<=2;bcd1<=6;bcd0<=3; end
			7264: begin bcd3<=7;bcd2<=2;bcd1<=6;bcd0<=4; end
			7265: begin bcd3<=7;bcd2<=2;bcd1<=6;bcd0<=5; end
			7266: begin bcd3<=7;bcd2<=2;bcd1<=6;bcd0<=6; end
			7267: begin bcd3<=7;bcd2<=2;bcd1<=6;bcd0<=7; end
			7268: begin bcd3<=7;bcd2<=2;bcd1<=6;bcd0<=8; end
			7269: begin bcd3<=7;bcd2<=2;bcd1<=6;bcd0<=9; end
			7270: begin bcd3<=7;bcd2<=2;bcd1<=7;bcd0<=0; end
			7271: begin bcd3<=7;bcd2<=2;bcd1<=7;bcd0<=1; end
			7272: begin bcd3<=7;bcd2<=2;bcd1<=7;bcd0<=2; end
			7273: begin bcd3<=7;bcd2<=2;bcd1<=7;bcd0<=3; end
			7274: begin bcd3<=7;bcd2<=2;bcd1<=7;bcd0<=4; end
			7275: begin bcd3<=7;bcd2<=2;bcd1<=7;bcd0<=5; end
			7276: begin bcd3<=7;bcd2<=2;bcd1<=7;bcd0<=6; end
			7277: begin bcd3<=7;bcd2<=2;bcd1<=7;bcd0<=7; end
			7278: begin bcd3<=7;bcd2<=2;bcd1<=7;bcd0<=8; end
			7279: begin bcd3<=7;bcd2<=2;bcd1<=7;bcd0<=9; end
			7280: begin bcd3<=7;bcd2<=2;bcd1<=8;bcd0<=0; end
			7281: begin bcd3<=7;bcd2<=2;bcd1<=8;bcd0<=1; end
			7282: begin bcd3<=7;bcd2<=2;bcd1<=8;bcd0<=2; end
			7283: begin bcd3<=7;bcd2<=2;bcd1<=8;bcd0<=3; end
			7284: begin bcd3<=7;bcd2<=2;bcd1<=8;bcd0<=4; end
			7285: begin bcd3<=7;bcd2<=2;bcd1<=8;bcd0<=5; end
			7286: begin bcd3<=7;bcd2<=2;bcd1<=8;bcd0<=6; end
			7287: begin bcd3<=7;bcd2<=2;bcd1<=8;bcd0<=7; end
			7288: begin bcd3<=7;bcd2<=2;bcd1<=8;bcd0<=8; end
			7289: begin bcd3<=7;bcd2<=2;bcd1<=8;bcd0<=9; end
			7290: begin bcd3<=7;bcd2<=2;bcd1<=9;bcd0<=0; end
			7291: begin bcd3<=7;bcd2<=2;bcd1<=9;bcd0<=1; end
			7292: begin bcd3<=7;bcd2<=2;bcd1<=9;bcd0<=2; end
			7293: begin bcd3<=7;bcd2<=2;bcd1<=9;bcd0<=3; end
			7294: begin bcd3<=7;bcd2<=2;bcd1<=9;bcd0<=4; end
			7295: begin bcd3<=7;bcd2<=2;bcd1<=9;bcd0<=5; end
			7296: begin bcd3<=7;bcd2<=2;bcd1<=9;bcd0<=6; end
			7297: begin bcd3<=7;bcd2<=2;bcd1<=9;bcd0<=7; end
			7298: begin bcd3<=7;bcd2<=2;bcd1<=9;bcd0<=8; end
			7299: begin bcd3<=7;bcd2<=2;bcd1<=9;bcd0<=9; end
			7300: begin bcd3<=7;bcd2<=3;bcd1<=0;bcd0<=0; end
			7301: begin bcd3<=7;bcd2<=3;bcd1<=0;bcd0<=1; end
			7302: begin bcd3<=7;bcd2<=3;bcd1<=0;bcd0<=2; end
			7303: begin bcd3<=7;bcd2<=3;bcd1<=0;bcd0<=3; end
			7304: begin bcd3<=7;bcd2<=3;bcd1<=0;bcd0<=4; end
			7305: begin bcd3<=7;bcd2<=3;bcd1<=0;bcd0<=5; end
			7306: begin bcd3<=7;bcd2<=3;bcd1<=0;bcd0<=6; end
			7307: begin bcd3<=7;bcd2<=3;bcd1<=0;bcd0<=7; end
			7308: begin bcd3<=7;bcd2<=3;bcd1<=0;bcd0<=8; end
			7309: begin bcd3<=7;bcd2<=3;bcd1<=0;bcd0<=9; end
			7310: begin bcd3<=7;bcd2<=3;bcd1<=1;bcd0<=0; end
			7311: begin bcd3<=7;bcd2<=3;bcd1<=1;bcd0<=1; end
			7312: begin bcd3<=7;bcd2<=3;bcd1<=1;bcd0<=2; end
			7313: begin bcd3<=7;bcd2<=3;bcd1<=1;bcd0<=3; end
			7314: begin bcd3<=7;bcd2<=3;bcd1<=1;bcd0<=4; end
			7315: begin bcd3<=7;bcd2<=3;bcd1<=1;bcd0<=5; end
			7316: begin bcd3<=7;bcd2<=3;bcd1<=1;bcd0<=6; end
			7317: begin bcd3<=7;bcd2<=3;bcd1<=1;bcd0<=7; end
			7318: begin bcd3<=7;bcd2<=3;bcd1<=1;bcd0<=8; end
			7319: begin bcd3<=7;bcd2<=3;bcd1<=1;bcd0<=9; end
			7320: begin bcd3<=7;bcd2<=3;bcd1<=2;bcd0<=0; end
			7321: begin bcd3<=7;bcd2<=3;bcd1<=2;bcd0<=1; end
			7322: begin bcd3<=7;bcd2<=3;bcd1<=2;bcd0<=2; end
			7323: begin bcd3<=7;bcd2<=3;bcd1<=2;bcd0<=3; end
			7324: begin bcd3<=7;bcd2<=3;bcd1<=2;bcd0<=4; end
			7325: begin bcd3<=7;bcd2<=3;bcd1<=2;bcd0<=5; end
			7326: begin bcd3<=7;bcd2<=3;bcd1<=2;bcd0<=6; end
			7327: begin bcd3<=7;bcd2<=3;bcd1<=2;bcd0<=7; end
			7328: begin bcd3<=7;bcd2<=3;bcd1<=2;bcd0<=8; end
			7329: begin bcd3<=7;bcd2<=3;bcd1<=2;bcd0<=9; end
			7330: begin bcd3<=7;bcd2<=3;bcd1<=3;bcd0<=0; end
			7331: begin bcd3<=7;bcd2<=3;bcd1<=3;bcd0<=1; end
			7332: begin bcd3<=7;bcd2<=3;bcd1<=3;bcd0<=2; end
			7333: begin bcd3<=7;bcd2<=3;bcd1<=3;bcd0<=3; end
			7334: begin bcd3<=7;bcd2<=3;bcd1<=3;bcd0<=4; end
			7335: begin bcd3<=7;bcd2<=3;bcd1<=3;bcd0<=5; end
			7336: begin bcd3<=7;bcd2<=3;bcd1<=3;bcd0<=6; end
			7337: begin bcd3<=7;bcd2<=3;bcd1<=3;bcd0<=7; end
			7338: begin bcd3<=7;bcd2<=3;bcd1<=3;bcd0<=8; end
			7339: begin bcd3<=7;bcd2<=3;bcd1<=3;bcd0<=9; end
			7340: begin bcd3<=7;bcd2<=3;bcd1<=4;bcd0<=0; end
			7341: begin bcd3<=7;bcd2<=3;bcd1<=4;bcd0<=1; end
			7342: begin bcd3<=7;bcd2<=3;bcd1<=4;bcd0<=2; end
			7343: begin bcd3<=7;bcd2<=3;bcd1<=4;bcd0<=3; end
			7344: begin bcd3<=7;bcd2<=3;bcd1<=4;bcd0<=4; end
			7345: begin bcd3<=7;bcd2<=3;bcd1<=4;bcd0<=5; end
			7346: begin bcd3<=7;bcd2<=3;bcd1<=4;bcd0<=6; end
			7347: begin bcd3<=7;bcd2<=3;bcd1<=4;bcd0<=7; end
			7348: begin bcd3<=7;bcd2<=3;bcd1<=4;bcd0<=8; end
			7349: begin bcd3<=7;bcd2<=3;bcd1<=4;bcd0<=9; end
			7350: begin bcd3<=7;bcd2<=3;bcd1<=5;bcd0<=0; end
			7351: begin bcd3<=7;bcd2<=3;bcd1<=5;bcd0<=1; end
			7352: begin bcd3<=7;bcd2<=3;bcd1<=5;bcd0<=2; end
			7353: begin bcd3<=7;bcd2<=3;bcd1<=5;bcd0<=3; end
			7354: begin bcd3<=7;bcd2<=3;bcd1<=5;bcd0<=4; end
			7355: begin bcd3<=7;bcd2<=3;bcd1<=5;bcd0<=5; end
			7356: begin bcd3<=7;bcd2<=3;bcd1<=5;bcd0<=6; end
			7357: begin bcd3<=7;bcd2<=3;bcd1<=5;bcd0<=7; end
			7358: begin bcd3<=7;bcd2<=3;bcd1<=5;bcd0<=8; end
			7359: begin bcd3<=7;bcd2<=3;bcd1<=5;bcd0<=9; end
			7360: begin bcd3<=7;bcd2<=3;bcd1<=6;bcd0<=0; end
			7361: begin bcd3<=7;bcd2<=3;bcd1<=6;bcd0<=1; end
			7362: begin bcd3<=7;bcd2<=3;bcd1<=6;bcd0<=2; end
			7363: begin bcd3<=7;bcd2<=3;bcd1<=6;bcd0<=3; end
			7364: begin bcd3<=7;bcd2<=3;bcd1<=6;bcd0<=4; end
			7365: begin bcd3<=7;bcd2<=3;bcd1<=6;bcd0<=5; end
			7366: begin bcd3<=7;bcd2<=3;bcd1<=6;bcd0<=6; end
			7367: begin bcd3<=7;bcd2<=3;bcd1<=6;bcd0<=7; end
			7368: begin bcd3<=7;bcd2<=3;bcd1<=6;bcd0<=8; end
			7369: begin bcd3<=7;bcd2<=3;bcd1<=6;bcd0<=9; end
			7370: begin bcd3<=7;bcd2<=3;bcd1<=7;bcd0<=0; end
			7371: begin bcd3<=7;bcd2<=3;bcd1<=7;bcd0<=1; end
			7372: begin bcd3<=7;bcd2<=3;bcd1<=7;bcd0<=2; end
			7373: begin bcd3<=7;bcd2<=3;bcd1<=7;bcd0<=3; end
			7374: begin bcd3<=7;bcd2<=3;bcd1<=7;bcd0<=4; end
			7375: begin bcd3<=7;bcd2<=3;bcd1<=7;bcd0<=5; end
			7376: begin bcd3<=7;bcd2<=3;bcd1<=7;bcd0<=6; end
			7377: begin bcd3<=7;bcd2<=3;bcd1<=7;bcd0<=7; end
			7378: begin bcd3<=7;bcd2<=3;bcd1<=7;bcd0<=8; end
			7379: begin bcd3<=7;bcd2<=3;bcd1<=7;bcd0<=9; end
			7380: begin bcd3<=7;bcd2<=3;bcd1<=8;bcd0<=0; end
			7381: begin bcd3<=7;bcd2<=3;bcd1<=8;bcd0<=1; end
			7382: begin bcd3<=7;bcd2<=3;bcd1<=8;bcd0<=2; end
			7383: begin bcd3<=7;bcd2<=3;bcd1<=8;bcd0<=3; end
			7384: begin bcd3<=7;bcd2<=3;bcd1<=8;bcd0<=4; end
			7385: begin bcd3<=7;bcd2<=3;bcd1<=8;bcd0<=5; end
			7386: begin bcd3<=7;bcd2<=3;bcd1<=8;bcd0<=6; end
			7387: begin bcd3<=7;bcd2<=3;bcd1<=8;bcd0<=7; end
			7388: begin bcd3<=7;bcd2<=3;bcd1<=8;bcd0<=8; end
			7389: begin bcd3<=7;bcd2<=3;bcd1<=8;bcd0<=9; end
			7390: begin bcd3<=7;bcd2<=3;bcd1<=9;bcd0<=0; end
			7391: begin bcd3<=7;bcd2<=3;bcd1<=9;bcd0<=1; end
			7392: begin bcd3<=7;bcd2<=3;bcd1<=9;bcd0<=2; end
			7393: begin bcd3<=7;bcd2<=3;bcd1<=9;bcd0<=3; end
			7394: begin bcd3<=7;bcd2<=3;bcd1<=9;bcd0<=4; end
			7395: begin bcd3<=7;bcd2<=3;bcd1<=9;bcd0<=5; end
			7396: begin bcd3<=7;bcd2<=3;bcd1<=9;bcd0<=6; end
			7397: begin bcd3<=7;bcd2<=3;bcd1<=9;bcd0<=7; end
			7398: begin bcd3<=7;bcd2<=3;bcd1<=9;bcd0<=8; end
			7399: begin bcd3<=7;bcd2<=3;bcd1<=9;bcd0<=9; end
			7400: begin bcd3<=7;bcd2<=4;bcd1<=0;bcd0<=0; end
			7401: begin bcd3<=7;bcd2<=4;bcd1<=0;bcd0<=1; end
			7402: begin bcd3<=7;bcd2<=4;bcd1<=0;bcd0<=2; end
			7403: begin bcd3<=7;bcd2<=4;bcd1<=0;bcd0<=3; end
			7404: begin bcd3<=7;bcd2<=4;bcd1<=0;bcd0<=4; end
			7405: begin bcd3<=7;bcd2<=4;bcd1<=0;bcd0<=5; end
			7406: begin bcd3<=7;bcd2<=4;bcd1<=0;bcd0<=6; end
			7407: begin bcd3<=7;bcd2<=4;bcd1<=0;bcd0<=7; end
			7408: begin bcd3<=7;bcd2<=4;bcd1<=0;bcd0<=8; end
			7409: begin bcd3<=7;bcd2<=4;bcd1<=0;bcd0<=9; end
			7410: begin bcd3<=7;bcd2<=4;bcd1<=1;bcd0<=0; end
			7411: begin bcd3<=7;bcd2<=4;bcd1<=1;bcd0<=1; end
			7412: begin bcd3<=7;bcd2<=4;bcd1<=1;bcd0<=2; end
			7413: begin bcd3<=7;bcd2<=4;bcd1<=1;bcd0<=3; end
			7414: begin bcd3<=7;bcd2<=4;bcd1<=1;bcd0<=4; end
			7415: begin bcd3<=7;bcd2<=4;bcd1<=1;bcd0<=5; end
			7416: begin bcd3<=7;bcd2<=4;bcd1<=1;bcd0<=6; end
			7417: begin bcd3<=7;bcd2<=4;bcd1<=1;bcd0<=7; end
			7418: begin bcd3<=7;bcd2<=4;bcd1<=1;bcd0<=8; end
			7419: begin bcd3<=7;bcd2<=4;bcd1<=1;bcd0<=9; end
			7420: begin bcd3<=7;bcd2<=4;bcd1<=2;bcd0<=0; end
			7421: begin bcd3<=7;bcd2<=4;bcd1<=2;bcd0<=1; end
			7422: begin bcd3<=7;bcd2<=4;bcd1<=2;bcd0<=2; end
			7423: begin bcd3<=7;bcd2<=4;bcd1<=2;bcd0<=3; end
			7424: begin bcd3<=7;bcd2<=4;bcd1<=2;bcd0<=4; end
			7425: begin bcd3<=7;bcd2<=4;bcd1<=2;bcd0<=5; end
			7426: begin bcd3<=7;bcd2<=4;bcd1<=2;bcd0<=6; end
			7427: begin bcd3<=7;bcd2<=4;bcd1<=2;bcd0<=7; end
			7428: begin bcd3<=7;bcd2<=4;bcd1<=2;bcd0<=8; end
			7429: begin bcd3<=7;bcd2<=4;bcd1<=2;bcd0<=9; end
			7430: begin bcd3<=7;bcd2<=4;bcd1<=3;bcd0<=0; end
			7431: begin bcd3<=7;bcd2<=4;bcd1<=3;bcd0<=1; end
			7432: begin bcd3<=7;bcd2<=4;bcd1<=3;bcd0<=2; end
			7433: begin bcd3<=7;bcd2<=4;bcd1<=3;bcd0<=3; end
			7434: begin bcd3<=7;bcd2<=4;bcd1<=3;bcd0<=4; end
			7435: begin bcd3<=7;bcd2<=4;bcd1<=3;bcd0<=5; end
			7436: begin bcd3<=7;bcd2<=4;bcd1<=3;bcd0<=6; end
			7437: begin bcd3<=7;bcd2<=4;bcd1<=3;bcd0<=7; end
			7438: begin bcd3<=7;bcd2<=4;bcd1<=3;bcd0<=8; end
			7439: begin bcd3<=7;bcd2<=4;bcd1<=3;bcd0<=9; end
			7440: begin bcd3<=7;bcd2<=4;bcd1<=4;bcd0<=0; end
			7441: begin bcd3<=7;bcd2<=4;bcd1<=4;bcd0<=1; end
			7442: begin bcd3<=7;bcd2<=4;bcd1<=4;bcd0<=2; end
			7443: begin bcd3<=7;bcd2<=4;bcd1<=4;bcd0<=3; end
			7444: begin bcd3<=7;bcd2<=4;bcd1<=4;bcd0<=4; end
			7445: begin bcd3<=7;bcd2<=4;bcd1<=4;bcd0<=5; end
			7446: begin bcd3<=7;bcd2<=4;bcd1<=4;bcd0<=6; end
			7447: begin bcd3<=7;bcd2<=4;bcd1<=4;bcd0<=7; end
			7448: begin bcd3<=7;bcd2<=4;bcd1<=4;bcd0<=8; end
			7449: begin bcd3<=7;bcd2<=4;bcd1<=4;bcd0<=9; end
			7450: begin bcd3<=7;bcd2<=4;bcd1<=5;bcd0<=0; end
			7451: begin bcd3<=7;bcd2<=4;bcd1<=5;bcd0<=1; end
			7452: begin bcd3<=7;bcd2<=4;bcd1<=5;bcd0<=2; end
			7453: begin bcd3<=7;bcd2<=4;bcd1<=5;bcd0<=3; end
			7454: begin bcd3<=7;bcd2<=4;bcd1<=5;bcd0<=4; end
			7455: begin bcd3<=7;bcd2<=4;bcd1<=5;bcd0<=5; end
			7456: begin bcd3<=7;bcd2<=4;bcd1<=5;bcd0<=6; end
			7457: begin bcd3<=7;bcd2<=4;bcd1<=5;bcd0<=7; end
			7458: begin bcd3<=7;bcd2<=4;bcd1<=5;bcd0<=8; end
			7459: begin bcd3<=7;bcd2<=4;bcd1<=5;bcd0<=9; end
			7460: begin bcd3<=7;bcd2<=4;bcd1<=6;bcd0<=0; end
			7461: begin bcd3<=7;bcd2<=4;bcd1<=6;bcd0<=1; end
			7462: begin bcd3<=7;bcd2<=4;bcd1<=6;bcd0<=2; end
			7463: begin bcd3<=7;bcd2<=4;bcd1<=6;bcd0<=3; end
			7464: begin bcd3<=7;bcd2<=4;bcd1<=6;bcd0<=4; end
			7465: begin bcd3<=7;bcd2<=4;bcd1<=6;bcd0<=5; end
			7466: begin bcd3<=7;bcd2<=4;bcd1<=6;bcd0<=6; end
			7467: begin bcd3<=7;bcd2<=4;bcd1<=6;bcd0<=7; end
			7468: begin bcd3<=7;bcd2<=4;bcd1<=6;bcd0<=8; end
			7469: begin bcd3<=7;bcd2<=4;bcd1<=6;bcd0<=9; end
			7470: begin bcd3<=7;bcd2<=4;bcd1<=7;bcd0<=0; end
			7471: begin bcd3<=7;bcd2<=4;bcd1<=7;bcd0<=1; end
			7472: begin bcd3<=7;bcd2<=4;bcd1<=7;bcd0<=2; end
			7473: begin bcd3<=7;bcd2<=4;bcd1<=7;bcd0<=3; end
			7474: begin bcd3<=7;bcd2<=4;bcd1<=7;bcd0<=4; end
			7475: begin bcd3<=7;bcd2<=4;bcd1<=7;bcd0<=5; end
			7476: begin bcd3<=7;bcd2<=4;bcd1<=7;bcd0<=6; end
			7477: begin bcd3<=7;bcd2<=4;bcd1<=7;bcd0<=7; end
			7478: begin bcd3<=7;bcd2<=4;bcd1<=7;bcd0<=8; end
			7479: begin bcd3<=7;bcd2<=4;bcd1<=7;bcd0<=9; end
			7480: begin bcd3<=7;bcd2<=4;bcd1<=8;bcd0<=0; end
			7481: begin bcd3<=7;bcd2<=4;bcd1<=8;bcd0<=1; end
			7482: begin bcd3<=7;bcd2<=4;bcd1<=8;bcd0<=2; end
			7483: begin bcd3<=7;bcd2<=4;bcd1<=8;bcd0<=3; end
			7484: begin bcd3<=7;bcd2<=4;bcd1<=8;bcd0<=4; end
			7485: begin bcd3<=7;bcd2<=4;bcd1<=8;bcd0<=5; end
			7486: begin bcd3<=7;bcd2<=4;bcd1<=8;bcd0<=6; end
			7487: begin bcd3<=7;bcd2<=4;bcd1<=8;bcd0<=7; end
			7488: begin bcd3<=7;bcd2<=4;bcd1<=8;bcd0<=8; end
			7489: begin bcd3<=7;bcd2<=4;bcd1<=8;bcd0<=9; end
			7490: begin bcd3<=7;bcd2<=4;bcd1<=9;bcd0<=0; end
			7491: begin bcd3<=7;bcd2<=4;bcd1<=9;bcd0<=1; end
			7492: begin bcd3<=7;bcd2<=4;bcd1<=9;bcd0<=2; end
			7493: begin bcd3<=7;bcd2<=4;bcd1<=9;bcd0<=3; end
			7494: begin bcd3<=7;bcd2<=4;bcd1<=9;bcd0<=4; end
			7495: begin bcd3<=7;bcd2<=4;bcd1<=9;bcd0<=5; end
			7496: begin bcd3<=7;bcd2<=4;bcd1<=9;bcd0<=6; end
			7497: begin bcd3<=7;bcd2<=4;bcd1<=9;bcd0<=7; end
			7498: begin bcd3<=7;bcd2<=4;bcd1<=9;bcd0<=8; end
			7499: begin bcd3<=7;bcd2<=4;bcd1<=9;bcd0<=9; end
			7500: begin bcd3<=7;bcd2<=5;bcd1<=0;bcd0<=0; end
			7501: begin bcd3<=7;bcd2<=5;bcd1<=0;bcd0<=1; end
			7502: begin bcd3<=7;bcd2<=5;bcd1<=0;bcd0<=2; end
			7503: begin bcd3<=7;bcd2<=5;bcd1<=0;bcd0<=3; end
			7504: begin bcd3<=7;bcd2<=5;bcd1<=0;bcd0<=4; end
			7505: begin bcd3<=7;bcd2<=5;bcd1<=0;bcd0<=5; end
			7506: begin bcd3<=7;bcd2<=5;bcd1<=0;bcd0<=6; end
			7507: begin bcd3<=7;bcd2<=5;bcd1<=0;bcd0<=7; end
			7508: begin bcd3<=7;bcd2<=5;bcd1<=0;bcd0<=8; end
			7509: begin bcd3<=7;bcd2<=5;bcd1<=0;bcd0<=9; end
			7510: begin bcd3<=7;bcd2<=5;bcd1<=1;bcd0<=0; end
			7511: begin bcd3<=7;bcd2<=5;bcd1<=1;bcd0<=1; end
			7512: begin bcd3<=7;bcd2<=5;bcd1<=1;bcd0<=2; end
			7513: begin bcd3<=7;bcd2<=5;bcd1<=1;bcd0<=3; end
			7514: begin bcd3<=7;bcd2<=5;bcd1<=1;bcd0<=4; end
			7515: begin bcd3<=7;bcd2<=5;bcd1<=1;bcd0<=5; end
			7516: begin bcd3<=7;bcd2<=5;bcd1<=1;bcd0<=6; end
			7517: begin bcd3<=7;bcd2<=5;bcd1<=1;bcd0<=7; end
			7518: begin bcd3<=7;bcd2<=5;bcd1<=1;bcd0<=8; end
			7519: begin bcd3<=7;bcd2<=5;bcd1<=1;bcd0<=9; end
			7520: begin bcd3<=7;bcd2<=5;bcd1<=2;bcd0<=0; end
			7521: begin bcd3<=7;bcd2<=5;bcd1<=2;bcd0<=1; end
			7522: begin bcd3<=7;bcd2<=5;bcd1<=2;bcd0<=2; end
			7523: begin bcd3<=7;bcd2<=5;bcd1<=2;bcd0<=3; end
			7524: begin bcd3<=7;bcd2<=5;bcd1<=2;bcd0<=4; end
			7525: begin bcd3<=7;bcd2<=5;bcd1<=2;bcd0<=5; end
			7526: begin bcd3<=7;bcd2<=5;bcd1<=2;bcd0<=6; end
			7527: begin bcd3<=7;bcd2<=5;bcd1<=2;bcd0<=7; end
			7528: begin bcd3<=7;bcd2<=5;bcd1<=2;bcd0<=8; end
			7529: begin bcd3<=7;bcd2<=5;bcd1<=2;bcd0<=9; end
			7530: begin bcd3<=7;bcd2<=5;bcd1<=3;bcd0<=0; end
			7531: begin bcd3<=7;bcd2<=5;bcd1<=3;bcd0<=1; end
			7532: begin bcd3<=7;bcd2<=5;bcd1<=3;bcd0<=2; end
			7533: begin bcd3<=7;bcd2<=5;bcd1<=3;bcd0<=3; end
			7534: begin bcd3<=7;bcd2<=5;bcd1<=3;bcd0<=4; end
			7535: begin bcd3<=7;bcd2<=5;bcd1<=3;bcd0<=5; end
			7536: begin bcd3<=7;bcd2<=5;bcd1<=3;bcd0<=6; end
			7537: begin bcd3<=7;bcd2<=5;bcd1<=3;bcd0<=7; end
			7538: begin bcd3<=7;bcd2<=5;bcd1<=3;bcd0<=8; end
			7539: begin bcd3<=7;bcd2<=5;bcd1<=3;bcd0<=9; end
			7540: begin bcd3<=7;bcd2<=5;bcd1<=4;bcd0<=0; end
			7541: begin bcd3<=7;bcd2<=5;bcd1<=4;bcd0<=1; end
			7542: begin bcd3<=7;bcd2<=5;bcd1<=4;bcd0<=2; end
			7543: begin bcd3<=7;bcd2<=5;bcd1<=4;bcd0<=3; end
			7544: begin bcd3<=7;bcd2<=5;bcd1<=4;bcd0<=4; end
			7545: begin bcd3<=7;bcd2<=5;bcd1<=4;bcd0<=5; end
			7546: begin bcd3<=7;bcd2<=5;bcd1<=4;bcd0<=6; end
			7547: begin bcd3<=7;bcd2<=5;bcd1<=4;bcd0<=7; end
			7548: begin bcd3<=7;bcd2<=5;bcd1<=4;bcd0<=8; end
			7549: begin bcd3<=7;bcd2<=5;bcd1<=4;bcd0<=9; end
			7550: begin bcd3<=7;bcd2<=5;bcd1<=5;bcd0<=0; end
			7551: begin bcd3<=7;bcd2<=5;bcd1<=5;bcd0<=1; end
			7552: begin bcd3<=7;bcd2<=5;bcd1<=5;bcd0<=2; end
			7553: begin bcd3<=7;bcd2<=5;bcd1<=5;bcd0<=3; end
			7554: begin bcd3<=7;bcd2<=5;bcd1<=5;bcd0<=4; end
			7555: begin bcd3<=7;bcd2<=5;bcd1<=5;bcd0<=5; end
			7556: begin bcd3<=7;bcd2<=5;bcd1<=5;bcd0<=6; end
			7557: begin bcd3<=7;bcd2<=5;bcd1<=5;bcd0<=7; end
			7558: begin bcd3<=7;bcd2<=5;bcd1<=5;bcd0<=8; end
			7559: begin bcd3<=7;bcd2<=5;bcd1<=5;bcd0<=9; end
			7560: begin bcd3<=7;bcd2<=5;bcd1<=6;bcd0<=0; end
			7561: begin bcd3<=7;bcd2<=5;bcd1<=6;bcd0<=1; end
			7562: begin bcd3<=7;bcd2<=5;bcd1<=6;bcd0<=2; end
			7563: begin bcd3<=7;bcd2<=5;bcd1<=6;bcd0<=3; end
			7564: begin bcd3<=7;bcd2<=5;bcd1<=6;bcd0<=4; end
			7565: begin bcd3<=7;bcd2<=5;bcd1<=6;bcd0<=5; end
			7566: begin bcd3<=7;bcd2<=5;bcd1<=6;bcd0<=6; end
			7567: begin bcd3<=7;bcd2<=5;bcd1<=6;bcd0<=7; end
			7568: begin bcd3<=7;bcd2<=5;bcd1<=6;bcd0<=8; end
			7569: begin bcd3<=7;bcd2<=5;bcd1<=6;bcd0<=9; end
			7570: begin bcd3<=7;bcd2<=5;bcd1<=7;bcd0<=0; end
			7571: begin bcd3<=7;bcd2<=5;bcd1<=7;bcd0<=1; end
			7572: begin bcd3<=7;bcd2<=5;bcd1<=7;bcd0<=2; end
			7573: begin bcd3<=7;bcd2<=5;bcd1<=7;bcd0<=3; end
			7574: begin bcd3<=7;bcd2<=5;bcd1<=7;bcd0<=4; end
			7575: begin bcd3<=7;bcd2<=5;bcd1<=7;bcd0<=5; end
			7576: begin bcd3<=7;bcd2<=5;bcd1<=7;bcd0<=6; end
			7577: begin bcd3<=7;bcd2<=5;bcd1<=7;bcd0<=7; end
			7578: begin bcd3<=7;bcd2<=5;bcd1<=7;bcd0<=8; end
			7579: begin bcd3<=7;bcd2<=5;bcd1<=7;bcd0<=9; end
			7580: begin bcd3<=7;bcd2<=5;bcd1<=8;bcd0<=0; end
			7581: begin bcd3<=7;bcd2<=5;bcd1<=8;bcd0<=1; end
			7582: begin bcd3<=7;bcd2<=5;bcd1<=8;bcd0<=2; end
			7583: begin bcd3<=7;bcd2<=5;bcd1<=8;bcd0<=3; end
			7584: begin bcd3<=7;bcd2<=5;bcd1<=8;bcd0<=4; end
			7585: begin bcd3<=7;bcd2<=5;bcd1<=8;bcd0<=5; end
			7586: begin bcd3<=7;bcd2<=5;bcd1<=8;bcd0<=6; end
			7587: begin bcd3<=7;bcd2<=5;bcd1<=8;bcd0<=7; end
			7588: begin bcd3<=7;bcd2<=5;bcd1<=8;bcd0<=8; end
			7589: begin bcd3<=7;bcd2<=5;bcd1<=8;bcd0<=9; end
			7590: begin bcd3<=7;bcd2<=5;bcd1<=9;bcd0<=0; end
			7591: begin bcd3<=7;bcd2<=5;bcd1<=9;bcd0<=1; end
			7592: begin bcd3<=7;bcd2<=5;bcd1<=9;bcd0<=2; end
			7593: begin bcd3<=7;bcd2<=5;bcd1<=9;bcd0<=3; end
			7594: begin bcd3<=7;bcd2<=5;bcd1<=9;bcd0<=4; end
			7595: begin bcd3<=7;bcd2<=5;bcd1<=9;bcd0<=5; end
			7596: begin bcd3<=7;bcd2<=5;bcd1<=9;bcd0<=6; end
			7597: begin bcd3<=7;bcd2<=5;bcd1<=9;bcd0<=7; end
			7598: begin bcd3<=7;bcd2<=5;bcd1<=9;bcd0<=8; end
			7599: begin bcd3<=7;bcd2<=5;bcd1<=9;bcd0<=9; end
			7600: begin bcd3<=7;bcd2<=6;bcd1<=0;bcd0<=0; end
			7601: begin bcd3<=7;bcd2<=6;bcd1<=0;bcd0<=1; end
			7602: begin bcd3<=7;bcd2<=6;bcd1<=0;bcd0<=2; end
			7603: begin bcd3<=7;bcd2<=6;bcd1<=0;bcd0<=3; end
			7604: begin bcd3<=7;bcd2<=6;bcd1<=0;bcd0<=4; end
			7605: begin bcd3<=7;bcd2<=6;bcd1<=0;bcd0<=5; end
			7606: begin bcd3<=7;bcd2<=6;bcd1<=0;bcd0<=6; end
			7607: begin bcd3<=7;bcd2<=6;bcd1<=0;bcd0<=7; end
			7608: begin bcd3<=7;bcd2<=6;bcd1<=0;bcd0<=8; end
			7609: begin bcd3<=7;bcd2<=6;bcd1<=0;bcd0<=9; end
			7610: begin bcd3<=7;bcd2<=6;bcd1<=1;bcd0<=0; end
			7611: begin bcd3<=7;bcd2<=6;bcd1<=1;bcd0<=1; end
			7612: begin bcd3<=7;bcd2<=6;bcd1<=1;bcd0<=2; end
			7613: begin bcd3<=7;bcd2<=6;bcd1<=1;bcd0<=3; end
			7614: begin bcd3<=7;bcd2<=6;bcd1<=1;bcd0<=4; end
			7615: begin bcd3<=7;bcd2<=6;bcd1<=1;bcd0<=5; end
			7616: begin bcd3<=7;bcd2<=6;bcd1<=1;bcd0<=6; end
			7617: begin bcd3<=7;bcd2<=6;bcd1<=1;bcd0<=7; end
			7618: begin bcd3<=7;bcd2<=6;bcd1<=1;bcd0<=8; end
			7619: begin bcd3<=7;bcd2<=6;bcd1<=1;bcd0<=9; end
			7620: begin bcd3<=7;bcd2<=6;bcd1<=2;bcd0<=0; end
			7621: begin bcd3<=7;bcd2<=6;bcd1<=2;bcd0<=1; end
			7622: begin bcd3<=7;bcd2<=6;bcd1<=2;bcd0<=2; end
			7623: begin bcd3<=7;bcd2<=6;bcd1<=2;bcd0<=3; end
			7624: begin bcd3<=7;bcd2<=6;bcd1<=2;bcd0<=4; end
			7625: begin bcd3<=7;bcd2<=6;bcd1<=2;bcd0<=5; end
			7626: begin bcd3<=7;bcd2<=6;bcd1<=2;bcd0<=6; end
			7627: begin bcd3<=7;bcd2<=6;bcd1<=2;bcd0<=7; end
			7628: begin bcd3<=7;bcd2<=6;bcd1<=2;bcd0<=8; end
			7629: begin bcd3<=7;bcd2<=6;bcd1<=2;bcd0<=9; end
			7630: begin bcd3<=7;bcd2<=6;bcd1<=3;bcd0<=0; end
			7631: begin bcd3<=7;bcd2<=6;bcd1<=3;bcd0<=1; end
			7632: begin bcd3<=7;bcd2<=6;bcd1<=3;bcd0<=2; end
			7633: begin bcd3<=7;bcd2<=6;bcd1<=3;bcd0<=3; end
			7634: begin bcd3<=7;bcd2<=6;bcd1<=3;bcd0<=4; end
			7635: begin bcd3<=7;bcd2<=6;bcd1<=3;bcd0<=5; end
			7636: begin bcd3<=7;bcd2<=6;bcd1<=3;bcd0<=6; end
			7637: begin bcd3<=7;bcd2<=6;bcd1<=3;bcd0<=7; end
			7638: begin bcd3<=7;bcd2<=6;bcd1<=3;bcd0<=8; end
			7639: begin bcd3<=7;bcd2<=6;bcd1<=3;bcd0<=9; end
			7640: begin bcd3<=7;bcd2<=6;bcd1<=4;bcd0<=0; end
			7641: begin bcd3<=7;bcd2<=6;bcd1<=4;bcd0<=1; end
			7642: begin bcd3<=7;bcd2<=6;bcd1<=4;bcd0<=2; end
			7643: begin bcd3<=7;bcd2<=6;bcd1<=4;bcd0<=3; end
			7644: begin bcd3<=7;bcd2<=6;bcd1<=4;bcd0<=4; end
			7645: begin bcd3<=7;bcd2<=6;bcd1<=4;bcd0<=5; end
			7646: begin bcd3<=7;bcd2<=6;bcd1<=4;bcd0<=6; end
			7647: begin bcd3<=7;bcd2<=6;bcd1<=4;bcd0<=7; end
			7648: begin bcd3<=7;bcd2<=6;bcd1<=4;bcd0<=8; end
			7649: begin bcd3<=7;bcd2<=6;bcd1<=4;bcd0<=9; end
			7650: begin bcd3<=7;bcd2<=6;bcd1<=5;bcd0<=0; end
			7651: begin bcd3<=7;bcd2<=6;bcd1<=5;bcd0<=1; end
			7652: begin bcd3<=7;bcd2<=6;bcd1<=5;bcd0<=2; end
			7653: begin bcd3<=7;bcd2<=6;bcd1<=5;bcd0<=3; end
			7654: begin bcd3<=7;bcd2<=6;bcd1<=5;bcd0<=4; end
			7655: begin bcd3<=7;bcd2<=6;bcd1<=5;bcd0<=5; end
			7656: begin bcd3<=7;bcd2<=6;bcd1<=5;bcd0<=6; end
			7657: begin bcd3<=7;bcd2<=6;bcd1<=5;bcd0<=7; end
			7658: begin bcd3<=7;bcd2<=6;bcd1<=5;bcd0<=8; end
			7659: begin bcd3<=7;bcd2<=6;bcd1<=5;bcd0<=9; end
			7660: begin bcd3<=7;bcd2<=6;bcd1<=6;bcd0<=0; end
			7661: begin bcd3<=7;bcd2<=6;bcd1<=6;bcd0<=1; end
			7662: begin bcd3<=7;bcd2<=6;bcd1<=6;bcd0<=2; end
			7663: begin bcd3<=7;bcd2<=6;bcd1<=6;bcd0<=3; end
			7664: begin bcd3<=7;bcd2<=6;bcd1<=6;bcd0<=4; end
			7665: begin bcd3<=7;bcd2<=6;bcd1<=6;bcd0<=5; end
			7666: begin bcd3<=7;bcd2<=6;bcd1<=6;bcd0<=6; end
			7667: begin bcd3<=7;bcd2<=6;bcd1<=6;bcd0<=7; end
			7668: begin bcd3<=7;bcd2<=6;bcd1<=6;bcd0<=8; end
			7669: begin bcd3<=7;bcd2<=6;bcd1<=6;bcd0<=9; end
			7670: begin bcd3<=7;bcd2<=6;bcd1<=7;bcd0<=0; end
			7671: begin bcd3<=7;bcd2<=6;bcd1<=7;bcd0<=1; end
			7672: begin bcd3<=7;bcd2<=6;bcd1<=7;bcd0<=2; end
			7673: begin bcd3<=7;bcd2<=6;bcd1<=7;bcd0<=3; end
			7674: begin bcd3<=7;bcd2<=6;bcd1<=7;bcd0<=4; end
			7675: begin bcd3<=7;bcd2<=6;bcd1<=7;bcd0<=5; end
			7676: begin bcd3<=7;bcd2<=6;bcd1<=7;bcd0<=6; end
			7677: begin bcd3<=7;bcd2<=6;bcd1<=7;bcd0<=7; end
			7678: begin bcd3<=7;bcd2<=6;bcd1<=7;bcd0<=8; end
			7679: begin bcd3<=7;bcd2<=6;bcd1<=7;bcd0<=9; end
			7680: begin bcd3<=7;bcd2<=6;bcd1<=8;bcd0<=0; end
			7681: begin bcd3<=7;bcd2<=6;bcd1<=8;bcd0<=1; end
			7682: begin bcd3<=7;bcd2<=6;bcd1<=8;bcd0<=2; end
			7683: begin bcd3<=7;bcd2<=6;bcd1<=8;bcd0<=3; end
			7684: begin bcd3<=7;bcd2<=6;bcd1<=8;bcd0<=4; end
			7685: begin bcd3<=7;bcd2<=6;bcd1<=8;bcd0<=5; end
			7686: begin bcd3<=7;bcd2<=6;bcd1<=8;bcd0<=6; end
			7687: begin bcd3<=7;bcd2<=6;bcd1<=8;bcd0<=7; end
			7688: begin bcd3<=7;bcd2<=6;bcd1<=8;bcd0<=8; end
			7689: begin bcd3<=7;bcd2<=6;bcd1<=8;bcd0<=9; end
			7690: begin bcd3<=7;bcd2<=6;bcd1<=9;bcd0<=0; end
			7691: begin bcd3<=7;bcd2<=6;bcd1<=9;bcd0<=1; end
			7692: begin bcd3<=7;bcd2<=6;bcd1<=9;bcd0<=2; end
			7693: begin bcd3<=7;bcd2<=6;bcd1<=9;bcd0<=3; end
			7694: begin bcd3<=7;bcd2<=6;bcd1<=9;bcd0<=4; end
			7695: begin bcd3<=7;bcd2<=6;bcd1<=9;bcd0<=5; end
			7696: begin bcd3<=7;bcd2<=6;bcd1<=9;bcd0<=6; end
			7697: begin bcd3<=7;bcd2<=6;bcd1<=9;bcd0<=7; end
			7698: begin bcd3<=7;bcd2<=6;bcd1<=9;bcd0<=8; end
			7699: begin bcd3<=7;bcd2<=6;bcd1<=9;bcd0<=9; end
			7700: begin bcd3<=7;bcd2<=7;bcd1<=0;bcd0<=0; end
			7701: begin bcd3<=7;bcd2<=7;bcd1<=0;bcd0<=1; end
			7702: begin bcd3<=7;bcd2<=7;bcd1<=0;bcd0<=2; end
			7703: begin bcd3<=7;bcd2<=7;bcd1<=0;bcd0<=3; end
			7704: begin bcd3<=7;bcd2<=7;bcd1<=0;bcd0<=4; end
			7705: begin bcd3<=7;bcd2<=7;bcd1<=0;bcd0<=5; end
			7706: begin bcd3<=7;bcd2<=7;bcd1<=0;bcd0<=6; end
			7707: begin bcd3<=7;bcd2<=7;bcd1<=0;bcd0<=7; end
			7708: begin bcd3<=7;bcd2<=7;bcd1<=0;bcd0<=8; end
			7709: begin bcd3<=7;bcd2<=7;bcd1<=0;bcd0<=9; end
			7710: begin bcd3<=7;bcd2<=7;bcd1<=1;bcd0<=0; end
			7711: begin bcd3<=7;bcd2<=7;bcd1<=1;bcd0<=1; end
			7712: begin bcd3<=7;bcd2<=7;bcd1<=1;bcd0<=2; end
			7713: begin bcd3<=7;bcd2<=7;bcd1<=1;bcd0<=3; end
			7714: begin bcd3<=7;bcd2<=7;bcd1<=1;bcd0<=4; end
			7715: begin bcd3<=7;bcd2<=7;bcd1<=1;bcd0<=5; end
			7716: begin bcd3<=7;bcd2<=7;bcd1<=1;bcd0<=6; end
			7717: begin bcd3<=7;bcd2<=7;bcd1<=1;bcd0<=7; end
			7718: begin bcd3<=7;bcd2<=7;bcd1<=1;bcd0<=8; end
			7719: begin bcd3<=7;bcd2<=7;bcd1<=1;bcd0<=9; end
			7720: begin bcd3<=7;bcd2<=7;bcd1<=2;bcd0<=0; end
			7721: begin bcd3<=7;bcd2<=7;bcd1<=2;bcd0<=1; end
			7722: begin bcd3<=7;bcd2<=7;bcd1<=2;bcd0<=2; end
			7723: begin bcd3<=7;bcd2<=7;bcd1<=2;bcd0<=3; end
			7724: begin bcd3<=7;bcd2<=7;bcd1<=2;bcd0<=4; end
			7725: begin bcd3<=7;bcd2<=7;bcd1<=2;bcd0<=5; end
			7726: begin bcd3<=7;bcd2<=7;bcd1<=2;bcd0<=6; end
			7727: begin bcd3<=7;bcd2<=7;bcd1<=2;bcd0<=7; end
			7728: begin bcd3<=7;bcd2<=7;bcd1<=2;bcd0<=8; end
			7729: begin bcd3<=7;bcd2<=7;bcd1<=2;bcd0<=9; end
			7730: begin bcd3<=7;bcd2<=7;bcd1<=3;bcd0<=0; end
			7731: begin bcd3<=7;bcd2<=7;bcd1<=3;bcd0<=1; end
			7732: begin bcd3<=7;bcd2<=7;bcd1<=3;bcd0<=2; end
			7733: begin bcd3<=7;bcd2<=7;bcd1<=3;bcd0<=3; end
			7734: begin bcd3<=7;bcd2<=7;bcd1<=3;bcd0<=4; end
			7735: begin bcd3<=7;bcd2<=7;bcd1<=3;bcd0<=5; end
			7736: begin bcd3<=7;bcd2<=7;bcd1<=3;bcd0<=6; end
			7737: begin bcd3<=7;bcd2<=7;bcd1<=3;bcd0<=7; end
			7738: begin bcd3<=7;bcd2<=7;bcd1<=3;bcd0<=8; end
			7739: begin bcd3<=7;bcd2<=7;bcd1<=3;bcd0<=9; end
			7740: begin bcd3<=7;bcd2<=7;bcd1<=4;bcd0<=0; end
			7741: begin bcd3<=7;bcd2<=7;bcd1<=4;bcd0<=1; end
			7742: begin bcd3<=7;bcd2<=7;bcd1<=4;bcd0<=2; end
			7743: begin bcd3<=7;bcd2<=7;bcd1<=4;bcd0<=3; end
			7744: begin bcd3<=7;bcd2<=7;bcd1<=4;bcd0<=4; end
			7745: begin bcd3<=7;bcd2<=7;bcd1<=4;bcd0<=5; end
			7746: begin bcd3<=7;bcd2<=7;bcd1<=4;bcd0<=6; end
			7747: begin bcd3<=7;bcd2<=7;bcd1<=4;bcd0<=7; end
			7748: begin bcd3<=7;bcd2<=7;bcd1<=4;bcd0<=8; end
			7749: begin bcd3<=7;bcd2<=7;bcd1<=4;bcd0<=9; end
			7750: begin bcd3<=7;bcd2<=7;bcd1<=5;bcd0<=0; end
			7751: begin bcd3<=7;bcd2<=7;bcd1<=5;bcd0<=1; end
			7752: begin bcd3<=7;bcd2<=7;bcd1<=5;bcd0<=2; end
			7753: begin bcd3<=7;bcd2<=7;bcd1<=5;bcd0<=3; end
			7754: begin bcd3<=7;bcd2<=7;bcd1<=5;bcd0<=4; end
			7755: begin bcd3<=7;bcd2<=7;bcd1<=5;bcd0<=5; end
			7756: begin bcd3<=7;bcd2<=7;bcd1<=5;bcd0<=6; end
			7757: begin bcd3<=7;bcd2<=7;bcd1<=5;bcd0<=7; end
			7758: begin bcd3<=7;bcd2<=7;bcd1<=5;bcd0<=8; end
			7759: begin bcd3<=7;bcd2<=7;bcd1<=5;bcd0<=9; end
			7760: begin bcd3<=7;bcd2<=7;bcd1<=6;bcd0<=0; end
			7761: begin bcd3<=7;bcd2<=7;bcd1<=6;bcd0<=1; end
			7762: begin bcd3<=7;bcd2<=7;bcd1<=6;bcd0<=2; end
			7763: begin bcd3<=7;bcd2<=7;bcd1<=6;bcd0<=3; end
			7764: begin bcd3<=7;bcd2<=7;bcd1<=6;bcd0<=4; end
			7765: begin bcd3<=7;bcd2<=7;bcd1<=6;bcd0<=5; end
			7766: begin bcd3<=7;bcd2<=7;bcd1<=6;bcd0<=6; end
			7767: begin bcd3<=7;bcd2<=7;bcd1<=6;bcd0<=7; end
			7768: begin bcd3<=7;bcd2<=7;bcd1<=6;bcd0<=8; end
			7769: begin bcd3<=7;bcd2<=7;bcd1<=6;bcd0<=9; end
			7770: begin bcd3<=7;bcd2<=7;bcd1<=7;bcd0<=0; end
			7771: begin bcd3<=7;bcd2<=7;bcd1<=7;bcd0<=1; end
			7772: begin bcd3<=7;bcd2<=7;bcd1<=7;bcd0<=2; end
			7773: begin bcd3<=7;bcd2<=7;bcd1<=7;bcd0<=3; end
			7774: begin bcd3<=7;bcd2<=7;bcd1<=7;bcd0<=4; end
			7775: begin bcd3<=7;bcd2<=7;bcd1<=7;bcd0<=5; end
			7776: begin bcd3<=7;bcd2<=7;bcd1<=7;bcd0<=6; end
			7777: begin bcd3<=7;bcd2<=7;bcd1<=7;bcd0<=7; end
			7778: begin bcd3<=7;bcd2<=7;bcd1<=7;bcd0<=8; end
			7779: begin bcd3<=7;bcd2<=7;bcd1<=7;bcd0<=9; end
			7780: begin bcd3<=7;bcd2<=7;bcd1<=8;bcd0<=0; end
			7781: begin bcd3<=7;bcd2<=7;bcd1<=8;bcd0<=1; end
			7782: begin bcd3<=7;bcd2<=7;bcd1<=8;bcd0<=2; end
			7783: begin bcd3<=7;bcd2<=7;bcd1<=8;bcd0<=3; end
			7784: begin bcd3<=7;bcd2<=7;bcd1<=8;bcd0<=4; end
			7785: begin bcd3<=7;bcd2<=7;bcd1<=8;bcd0<=5; end
			7786: begin bcd3<=7;bcd2<=7;bcd1<=8;bcd0<=6; end
			7787: begin bcd3<=7;bcd2<=7;bcd1<=8;bcd0<=7; end
			7788: begin bcd3<=7;bcd2<=7;bcd1<=8;bcd0<=8; end
			7789: begin bcd3<=7;bcd2<=7;bcd1<=8;bcd0<=9; end
			7790: begin bcd3<=7;bcd2<=7;bcd1<=9;bcd0<=0; end
			7791: begin bcd3<=7;bcd2<=7;bcd1<=9;bcd0<=1; end
			7792: begin bcd3<=7;bcd2<=7;bcd1<=9;bcd0<=2; end
			7793: begin bcd3<=7;bcd2<=7;bcd1<=9;bcd0<=3; end
			7794: begin bcd3<=7;bcd2<=7;bcd1<=9;bcd0<=4; end
			7795: begin bcd3<=7;bcd2<=7;bcd1<=9;bcd0<=5; end
			7796: begin bcd3<=7;bcd2<=7;bcd1<=9;bcd0<=6; end
			7797: begin bcd3<=7;bcd2<=7;bcd1<=9;bcd0<=7; end
			7798: begin bcd3<=7;bcd2<=7;bcd1<=9;bcd0<=8; end
			7799: begin bcd3<=7;bcd2<=7;bcd1<=9;bcd0<=9; end
			7800: begin bcd3<=7;bcd2<=8;bcd1<=0;bcd0<=0; end
			7801: begin bcd3<=7;bcd2<=8;bcd1<=0;bcd0<=1; end
			7802: begin bcd3<=7;bcd2<=8;bcd1<=0;bcd0<=2; end
			7803: begin bcd3<=7;bcd2<=8;bcd1<=0;bcd0<=3; end
			7804: begin bcd3<=7;bcd2<=8;bcd1<=0;bcd0<=4; end
			7805: begin bcd3<=7;bcd2<=8;bcd1<=0;bcd0<=5; end
			7806: begin bcd3<=7;bcd2<=8;bcd1<=0;bcd0<=6; end
			7807: begin bcd3<=7;bcd2<=8;bcd1<=0;bcd0<=7; end
			7808: begin bcd3<=7;bcd2<=8;bcd1<=0;bcd0<=8; end
			7809: begin bcd3<=7;bcd2<=8;bcd1<=0;bcd0<=9; end
			7810: begin bcd3<=7;bcd2<=8;bcd1<=1;bcd0<=0; end
			7811: begin bcd3<=7;bcd2<=8;bcd1<=1;bcd0<=1; end
			7812: begin bcd3<=7;bcd2<=8;bcd1<=1;bcd0<=2; end
			7813: begin bcd3<=7;bcd2<=8;bcd1<=1;bcd0<=3; end
			7814: begin bcd3<=7;bcd2<=8;bcd1<=1;bcd0<=4; end
			7815: begin bcd3<=7;bcd2<=8;bcd1<=1;bcd0<=5; end
			7816: begin bcd3<=7;bcd2<=8;bcd1<=1;bcd0<=6; end
			7817: begin bcd3<=7;bcd2<=8;bcd1<=1;bcd0<=7; end
			7818: begin bcd3<=7;bcd2<=8;bcd1<=1;bcd0<=8; end
			7819: begin bcd3<=7;bcd2<=8;bcd1<=1;bcd0<=9; end
			7820: begin bcd3<=7;bcd2<=8;bcd1<=2;bcd0<=0; end
			7821: begin bcd3<=7;bcd2<=8;bcd1<=2;bcd0<=1; end
			7822: begin bcd3<=7;bcd2<=8;bcd1<=2;bcd0<=2; end
			7823: begin bcd3<=7;bcd2<=8;bcd1<=2;bcd0<=3; end
			7824: begin bcd3<=7;bcd2<=8;bcd1<=2;bcd0<=4; end
			7825: begin bcd3<=7;bcd2<=8;bcd1<=2;bcd0<=5; end
			7826: begin bcd3<=7;bcd2<=8;bcd1<=2;bcd0<=6; end
			7827: begin bcd3<=7;bcd2<=8;bcd1<=2;bcd0<=7; end
			7828: begin bcd3<=7;bcd2<=8;bcd1<=2;bcd0<=8; end
			7829: begin bcd3<=7;bcd2<=8;bcd1<=2;bcd0<=9; end
			7830: begin bcd3<=7;bcd2<=8;bcd1<=3;bcd0<=0; end
			7831: begin bcd3<=7;bcd2<=8;bcd1<=3;bcd0<=1; end
			7832: begin bcd3<=7;bcd2<=8;bcd1<=3;bcd0<=2; end
			7833: begin bcd3<=7;bcd2<=8;bcd1<=3;bcd0<=3; end
			7834: begin bcd3<=7;bcd2<=8;bcd1<=3;bcd0<=4; end
			7835: begin bcd3<=7;bcd2<=8;bcd1<=3;bcd0<=5; end
			7836: begin bcd3<=7;bcd2<=8;bcd1<=3;bcd0<=6; end
			7837: begin bcd3<=7;bcd2<=8;bcd1<=3;bcd0<=7; end
			7838: begin bcd3<=7;bcd2<=8;bcd1<=3;bcd0<=8; end
			7839: begin bcd3<=7;bcd2<=8;bcd1<=3;bcd0<=9; end
			7840: begin bcd3<=7;bcd2<=8;bcd1<=4;bcd0<=0; end
			7841: begin bcd3<=7;bcd2<=8;bcd1<=4;bcd0<=1; end
			7842: begin bcd3<=7;bcd2<=8;bcd1<=4;bcd0<=2; end
			7843: begin bcd3<=7;bcd2<=8;bcd1<=4;bcd0<=3; end
			7844: begin bcd3<=7;bcd2<=8;bcd1<=4;bcd0<=4; end
			7845: begin bcd3<=7;bcd2<=8;bcd1<=4;bcd0<=5; end
			7846: begin bcd3<=7;bcd2<=8;bcd1<=4;bcd0<=6; end
			7847: begin bcd3<=7;bcd2<=8;bcd1<=4;bcd0<=7; end
			7848: begin bcd3<=7;bcd2<=8;bcd1<=4;bcd0<=8; end
			7849: begin bcd3<=7;bcd2<=8;bcd1<=4;bcd0<=9; end
			7850: begin bcd3<=7;bcd2<=8;bcd1<=5;bcd0<=0; end
			7851: begin bcd3<=7;bcd2<=8;bcd1<=5;bcd0<=1; end
			7852: begin bcd3<=7;bcd2<=8;bcd1<=5;bcd0<=2; end
			7853: begin bcd3<=7;bcd2<=8;bcd1<=5;bcd0<=3; end
			7854: begin bcd3<=7;bcd2<=8;bcd1<=5;bcd0<=4; end
			7855: begin bcd3<=7;bcd2<=8;bcd1<=5;bcd0<=5; end
			7856: begin bcd3<=7;bcd2<=8;bcd1<=5;bcd0<=6; end
			7857: begin bcd3<=7;bcd2<=8;bcd1<=5;bcd0<=7; end
			7858: begin bcd3<=7;bcd2<=8;bcd1<=5;bcd0<=8; end
			7859: begin bcd3<=7;bcd2<=8;bcd1<=5;bcd0<=9; end
			7860: begin bcd3<=7;bcd2<=8;bcd1<=6;bcd0<=0; end
			7861: begin bcd3<=7;bcd2<=8;bcd1<=6;bcd0<=1; end
			7862: begin bcd3<=7;bcd2<=8;bcd1<=6;bcd0<=2; end
			7863: begin bcd3<=7;bcd2<=8;bcd1<=6;bcd0<=3; end
			7864: begin bcd3<=7;bcd2<=8;bcd1<=6;bcd0<=4; end
			7865: begin bcd3<=7;bcd2<=8;bcd1<=6;bcd0<=5; end
			7866: begin bcd3<=7;bcd2<=8;bcd1<=6;bcd0<=6; end
			7867: begin bcd3<=7;bcd2<=8;bcd1<=6;bcd0<=7; end
			7868: begin bcd3<=7;bcd2<=8;bcd1<=6;bcd0<=8; end
			7869: begin bcd3<=7;bcd2<=8;bcd1<=6;bcd0<=9; end
			7870: begin bcd3<=7;bcd2<=8;bcd1<=7;bcd0<=0; end
			7871: begin bcd3<=7;bcd2<=8;bcd1<=7;bcd0<=1; end
			7872: begin bcd3<=7;bcd2<=8;bcd1<=7;bcd0<=2; end
			7873: begin bcd3<=7;bcd2<=8;bcd1<=7;bcd0<=3; end
			7874: begin bcd3<=7;bcd2<=8;bcd1<=7;bcd0<=4; end
			7875: begin bcd3<=7;bcd2<=8;bcd1<=7;bcd0<=5; end
			7876: begin bcd3<=7;bcd2<=8;bcd1<=7;bcd0<=6; end
			7877: begin bcd3<=7;bcd2<=8;bcd1<=7;bcd0<=7; end
			7878: begin bcd3<=7;bcd2<=8;bcd1<=7;bcd0<=8; end
			7879: begin bcd3<=7;bcd2<=8;bcd1<=7;bcd0<=9; end
			7880: begin bcd3<=7;bcd2<=8;bcd1<=8;bcd0<=0; end
			7881: begin bcd3<=7;bcd2<=8;bcd1<=8;bcd0<=1; end
			7882: begin bcd3<=7;bcd2<=8;bcd1<=8;bcd0<=2; end
			7883: begin bcd3<=7;bcd2<=8;bcd1<=8;bcd0<=3; end
			7884: begin bcd3<=7;bcd2<=8;bcd1<=8;bcd0<=4; end
			7885: begin bcd3<=7;bcd2<=8;bcd1<=8;bcd0<=5; end
			7886: begin bcd3<=7;bcd2<=8;bcd1<=8;bcd0<=6; end
			7887: begin bcd3<=7;bcd2<=8;bcd1<=8;bcd0<=7; end
			7888: begin bcd3<=7;bcd2<=8;bcd1<=8;bcd0<=8; end
			7889: begin bcd3<=7;bcd2<=8;bcd1<=8;bcd0<=9; end
			7890: begin bcd3<=7;bcd2<=8;bcd1<=9;bcd0<=0; end
			7891: begin bcd3<=7;bcd2<=8;bcd1<=9;bcd0<=1; end
			7892: begin bcd3<=7;bcd2<=8;bcd1<=9;bcd0<=2; end
			7893: begin bcd3<=7;bcd2<=8;bcd1<=9;bcd0<=3; end
			7894: begin bcd3<=7;bcd2<=8;bcd1<=9;bcd0<=4; end
			7895: begin bcd3<=7;bcd2<=8;bcd1<=9;bcd0<=5; end
			7896: begin bcd3<=7;bcd2<=8;bcd1<=9;bcd0<=6; end
			7897: begin bcd3<=7;bcd2<=8;bcd1<=9;bcd0<=7; end
			7898: begin bcd3<=7;bcd2<=8;bcd1<=9;bcd0<=8; end
			7899: begin bcd3<=7;bcd2<=8;bcd1<=9;bcd0<=9; end
			7900: begin bcd3<=7;bcd2<=9;bcd1<=0;bcd0<=0; end
			7901: begin bcd3<=7;bcd2<=9;bcd1<=0;bcd0<=1; end
			7902: begin bcd3<=7;bcd2<=9;bcd1<=0;bcd0<=2; end
			7903: begin bcd3<=7;bcd2<=9;bcd1<=0;bcd0<=3; end
			7904: begin bcd3<=7;bcd2<=9;bcd1<=0;bcd0<=4; end
			7905: begin bcd3<=7;bcd2<=9;bcd1<=0;bcd0<=5; end
			7906: begin bcd3<=7;bcd2<=9;bcd1<=0;bcd0<=6; end
			7907: begin bcd3<=7;bcd2<=9;bcd1<=0;bcd0<=7; end
			7908: begin bcd3<=7;bcd2<=9;bcd1<=0;bcd0<=8; end
			7909: begin bcd3<=7;bcd2<=9;bcd1<=0;bcd0<=9; end
			7910: begin bcd3<=7;bcd2<=9;bcd1<=1;bcd0<=0; end
			7911: begin bcd3<=7;bcd2<=9;bcd1<=1;bcd0<=1; end
			7912: begin bcd3<=7;bcd2<=9;bcd1<=1;bcd0<=2; end
			7913: begin bcd3<=7;bcd2<=9;bcd1<=1;bcd0<=3; end
			7914: begin bcd3<=7;bcd2<=9;bcd1<=1;bcd0<=4; end
			7915: begin bcd3<=7;bcd2<=9;bcd1<=1;bcd0<=5; end
			7916: begin bcd3<=7;bcd2<=9;bcd1<=1;bcd0<=6; end
			7917: begin bcd3<=7;bcd2<=9;bcd1<=1;bcd0<=7; end
			7918: begin bcd3<=7;bcd2<=9;bcd1<=1;bcd0<=8; end
			7919: begin bcd3<=7;bcd2<=9;bcd1<=1;bcd0<=9; end
			7920: begin bcd3<=7;bcd2<=9;bcd1<=2;bcd0<=0; end
			7921: begin bcd3<=7;bcd2<=9;bcd1<=2;bcd0<=1; end
			7922: begin bcd3<=7;bcd2<=9;bcd1<=2;bcd0<=2; end
			7923: begin bcd3<=7;bcd2<=9;bcd1<=2;bcd0<=3; end
			7924: begin bcd3<=7;bcd2<=9;bcd1<=2;bcd0<=4; end
			7925: begin bcd3<=7;bcd2<=9;bcd1<=2;bcd0<=5; end
			7926: begin bcd3<=7;bcd2<=9;bcd1<=2;bcd0<=6; end
			7927: begin bcd3<=7;bcd2<=9;bcd1<=2;bcd0<=7; end
			7928: begin bcd3<=7;bcd2<=9;bcd1<=2;bcd0<=8; end
			7929: begin bcd3<=7;bcd2<=9;bcd1<=2;bcd0<=9; end
			7930: begin bcd3<=7;bcd2<=9;bcd1<=3;bcd0<=0; end
			7931: begin bcd3<=7;bcd2<=9;bcd1<=3;bcd0<=1; end
			7932: begin bcd3<=7;bcd2<=9;bcd1<=3;bcd0<=2; end
			7933: begin bcd3<=7;bcd2<=9;bcd1<=3;bcd0<=3; end
			7934: begin bcd3<=7;bcd2<=9;bcd1<=3;bcd0<=4; end
			7935: begin bcd3<=7;bcd2<=9;bcd1<=3;bcd0<=5; end
			7936: begin bcd3<=7;bcd2<=9;bcd1<=3;bcd0<=6; end
			7937: begin bcd3<=7;bcd2<=9;bcd1<=3;bcd0<=7; end
			7938: begin bcd3<=7;bcd2<=9;bcd1<=3;bcd0<=8; end
			7939: begin bcd3<=7;bcd2<=9;bcd1<=3;bcd0<=9; end
			7940: begin bcd3<=7;bcd2<=9;bcd1<=4;bcd0<=0; end
			7941: begin bcd3<=7;bcd2<=9;bcd1<=4;bcd0<=1; end
			7942: begin bcd3<=7;bcd2<=9;bcd1<=4;bcd0<=2; end
			7943: begin bcd3<=7;bcd2<=9;bcd1<=4;bcd0<=3; end
			7944: begin bcd3<=7;bcd2<=9;bcd1<=4;bcd0<=4; end
			7945: begin bcd3<=7;bcd2<=9;bcd1<=4;bcd0<=5; end
			7946: begin bcd3<=7;bcd2<=9;bcd1<=4;bcd0<=6; end
			7947: begin bcd3<=7;bcd2<=9;bcd1<=4;bcd0<=7; end
			7948: begin bcd3<=7;bcd2<=9;bcd1<=4;bcd0<=8; end
			7949: begin bcd3<=7;bcd2<=9;bcd1<=4;bcd0<=9; end
			7950: begin bcd3<=7;bcd2<=9;bcd1<=5;bcd0<=0; end
			7951: begin bcd3<=7;bcd2<=9;bcd1<=5;bcd0<=1; end
			7952: begin bcd3<=7;bcd2<=9;bcd1<=5;bcd0<=2; end
			7953: begin bcd3<=7;bcd2<=9;bcd1<=5;bcd0<=3; end
			7954: begin bcd3<=7;bcd2<=9;bcd1<=5;bcd0<=4; end
			7955: begin bcd3<=7;bcd2<=9;bcd1<=5;bcd0<=5; end
			7956: begin bcd3<=7;bcd2<=9;bcd1<=5;bcd0<=6; end
			7957: begin bcd3<=7;bcd2<=9;bcd1<=5;bcd0<=7; end
			7958: begin bcd3<=7;bcd2<=9;bcd1<=5;bcd0<=8; end
			7959: begin bcd3<=7;bcd2<=9;bcd1<=5;bcd0<=9; end
			7960: begin bcd3<=7;bcd2<=9;bcd1<=6;bcd0<=0; end
			7961: begin bcd3<=7;bcd2<=9;bcd1<=6;bcd0<=1; end
			7962: begin bcd3<=7;bcd2<=9;bcd1<=6;bcd0<=2; end
			7963: begin bcd3<=7;bcd2<=9;bcd1<=6;bcd0<=3; end
			7964: begin bcd3<=7;bcd2<=9;bcd1<=6;bcd0<=4; end
			7965: begin bcd3<=7;bcd2<=9;bcd1<=6;bcd0<=5; end
			7966: begin bcd3<=7;bcd2<=9;bcd1<=6;bcd0<=6; end
			7967: begin bcd3<=7;bcd2<=9;bcd1<=6;bcd0<=7; end
			7968: begin bcd3<=7;bcd2<=9;bcd1<=6;bcd0<=8; end
			7969: begin bcd3<=7;bcd2<=9;bcd1<=6;bcd0<=9; end
			7970: begin bcd3<=7;bcd2<=9;bcd1<=7;bcd0<=0; end
			7971: begin bcd3<=7;bcd2<=9;bcd1<=7;bcd0<=1; end
			7972: begin bcd3<=7;bcd2<=9;bcd1<=7;bcd0<=2; end
			7973: begin bcd3<=7;bcd2<=9;bcd1<=7;bcd0<=3; end
			7974: begin bcd3<=7;bcd2<=9;bcd1<=7;bcd0<=4; end
			7975: begin bcd3<=7;bcd2<=9;bcd1<=7;bcd0<=5; end
			7976: begin bcd3<=7;bcd2<=9;bcd1<=7;bcd0<=6; end
			7977: begin bcd3<=7;bcd2<=9;bcd1<=7;bcd0<=7; end
			7978: begin bcd3<=7;bcd2<=9;bcd1<=7;bcd0<=8; end
			7979: begin bcd3<=7;bcd2<=9;bcd1<=7;bcd0<=9; end
			7980: begin bcd3<=7;bcd2<=9;bcd1<=8;bcd0<=0; end
			7981: begin bcd3<=7;bcd2<=9;bcd1<=8;bcd0<=1; end
			7982: begin bcd3<=7;bcd2<=9;bcd1<=8;bcd0<=2; end
			7983: begin bcd3<=7;bcd2<=9;bcd1<=8;bcd0<=3; end
			7984: begin bcd3<=7;bcd2<=9;bcd1<=8;bcd0<=4; end
			7985: begin bcd3<=7;bcd2<=9;bcd1<=8;bcd0<=5; end
			7986: begin bcd3<=7;bcd2<=9;bcd1<=8;bcd0<=6; end
			7987: begin bcd3<=7;bcd2<=9;bcd1<=8;bcd0<=7; end
			7988: begin bcd3<=7;bcd2<=9;bcd1<=8;bcd0<=8; end
			7989: begin bcd3<=7;bcd2<=9;bcd1<=8;bcd0<=9; end
			7990: begin bcd3<=7;bcd2<=9;bcd1<=9;bcd0<=0; end
			7991: begin bcd3<=7;bcd2<=9;bcd1<=9;bcd0<=1; end
			7992: begin bcd3<=7;bcd2<=9;bcd1<=9;bcd0<=2; end
			7993: begin bcd3<=7;bcd2<=9;bcd1<=9;bcd0<=3; end
			7994: begin bcd3<=7;bcd2<=9;bcd1<=9;bcd0<=4; end
			7995: begin bcd3<=7;bcd2<=9;bcd1<=9;bcd0<=5; end
			7996: begin bcd3<=7;bcd2<=9;bcd1<=9;bcd0<=6; end
			7997: begin bcd3<=7;bcd2<=9;bcd1<=9;bcd0<=7; end
			7998: begin bcd3<=7;bcd2<=9;bcd1<=9;bcd0<=8; end
			7999: begin bcd3<=7;bcd2<=9;bcd1<=9;bcd0<=9; end
			8000: begin bcd3<=8;bcd2<=0;bcd1<=0;bcd0<=0; end
			8001: begin bcd3<=8;bcd2<=0;bcd1<=0;bcd0<=1; end
			8002: begin bcd3<=8;bcd2<=0;bcd1<=0;bcd0<=2; end
			8003: begin bcd3<=8;bcd2<=0;bcd1<=0;bcd0<=3; end
			8004: begin bcd3<=8;bcd2<=0;bcd1<=0;bcd0<=4; end
			8005: begin bcd3<=8;bcd2<=0;bcd1<=0;bcd0<=5; end
			8006: begin bcd3<=8;bcd2<=0;bcd1<=0;bcd0<=6; end
			8007: begin bcd3<=8;bcd2<=0;bcd1<=0;bcd0<=7; end
			8008: begin bcd3<=8;bcd2<=0;bcd1<=0;bcd0<=8; end
			8009: begin bcd3<=8;bcd2<=0;bcd1<=0;bcd0<=9; end
			8010: begin bcd3<=8;bcd2<=0;bcd1<=1;bcd0<=0; end
			8011: begin bcd3<=8;bcd2<=0;bcd1<=1;bcd0<=1; end
			8012: begin bcd3<=8;bcd2<=0;bcd1<=1;bcd0<=2; end
			8013: begin bcd3<=8;bcd2<=0;bcd1<=1;bcd0<=3; end
			8014: begin bcd3<=8;bcd2<=0;bcd1<=1;bcd0<=4; end
			8015: begin bcd3<=8;bcd2<=0;bcd1<=1;bcd0<=5; end
			8016: begin bcd3<=8;bcd2<=0;bcd1<=1;bcd0<=6; end
			8017: begin bcd3<=8;bcd2<=0;bcd1<=1;bcd0<=7; end
			8018: begin bcd3<=8;bcd2<=0;bcd1<=1;bcd0<=8; end
			8019: begin bcd3<=8;bcd2<=0;bcd1<=1;bcd0<=9; end
			8020: begin bcd3<=8;bcd2<=0;bcd1<=2;bcd0<=0; end
			8021: begin bcd3<=8;bcd2<=0;bcd1<=2;bcd0<=1; end
			8022: begin bcd3<=8;bcd2<=0;bcd1<=2;bcd0<=2; end
			8023: begin bcd3<=8;bcd2<=0;bcd1<=2;bcd0<=3; end
			8024: begin bcd3<=8;bcd2<=0;bcd1<=2;bcd0<=4; end
			8025: begin bcd3<=8;bcd2<=0;bcd1<=2;bcd0<=5; end
			8026: begin bcd3<=8;bcd2<=0;bcd1<=2;bcd0<=6; end
			8027: begin bcd3<=8;bcd2<=0;bcd1<=2;bcd0<=7; end
			8028: begin bcd3<=8;bcd2<=0;bcd1<=2;bcd0<=8; end
			8029: begin bcd3<=8;bcd2<=0;bcd1<=2;bcd0<=9; end
			8030: begin bcd3<=8;bcd2<=0;bcd1<=3;bcd0<=0; end
			8031: begin bcd3<=8;bcd2<=0;bcd1<=3;bcd0<=1; end
			8032: begin bcd3<=8;bcd2<=0;bcd1<=3;bcd0<=2; end
			8033: begin bcd3<=8;bcd2<=0;bcd1<=3;bcd0<=3; end
			8034: begin bcd3<=8;bcd2<=0;bcd1<=3;bcd0<=4; end
			8035: begin bcd3<=8;bcd2<=0;bcd1<=3;bcd0<=5; end
			8036: begin bcd3<=8;bcd2<=0;bcd1<=3;bcd0<=6; end
			8037: begin bcd3<=8;bcd2<=0;bcd1<=3;bcd0<=7; end
			8038: begin bcd3<=8;bcd2<=0;bcd1<=3;bcd0<=8; end
			8039: begin bcd3<=8;bcd2<=0;bcd1<=3;bcd0<=9; end
			8040: begin bcd3<=8;bcd2<=0;bcd1<=4;bcd0<=0; end
			8041: begin bcd3<=8;bcd2<=0;bcd1<=4;bcd0<=1; end
			8042: begin bcd3<=8;bcd2<=0;bcd1<=4;bcd0<=2; end
			8043: begin bcd3<=8;bcd2<=0;bcd1<=4;bcd0<=3; end
			8044: begin bcd3<=8;bcd2<=0;bcd1<=4;bcd0<=4; end
			8045: begin bcd3<=8;bcd2<=0;bcd1<=4;bcd0<=5; end
			8046: begin bcd3<=8;bcd2<=0;bcd1<=4;bcd0<=6; end
			8047: begin bcd3<=8;bcd2<=0;bcd1<=4;bcd0<=7; end
			8048: begin bcd3<=8;bcd2<=0;bcd1<=4;bcd0<=8; end
			8049: begin bcd3<=8;bcd2<=0;bcd1<=4;bcd0<=9; end
			8050: begin bcd3<=8;bcd2<=0;bcd1<=5;bcd0<=0; end
			8051: begin bcd3<=8;bcd2<=0;bcd1<=5;bcd0<=1; end
			8052: begin bcd3<=8;bcd2<=0;bcd1<=5;bcd0<=2; end
			8053: begin bcd3<=8;bcd2<=0;bcd1<=5;bcd0<=3; end
			8054: begin bcd3<=8;bcd2<=0;bcd1<=5;bcd0<=4; end
			8055: begin bcd3<=8;bcd2<=0;bcd1<=5;bcd0<=5; end
			8056: begin bcd3<=8;bcd2<=0;bcd1<=5;bcd0<=6; end
			8057: begin bcd3<=8;bcd2<=0;bcd1<=5;bcd0<=7; end
			8058: begin bcd3<=8;bcd2<=0;bcd1<=5;bcd0<=8; end
			8059: begin bcd3<=8;bcd2<=0;bcd1<=5;bcd0<=9; end
			8060: begin bcd3<=8;bcd2<=0;bcd1<=6;bcd0<=0; end
			8061: begin bcd3<=8;bcd2<=0;bcd1<=6;bcd0<=1; end
			8062: begin bcd3<=8;bcd2<=0;bcd1<=6;bcd0<=2; end
			8063: begin bcd3<=8;bcd2<=0;bcd1<=6;bcd0<=3; end
			8064: begin bcd3<=8;bcd2<=0;bcd1<=6;bcd0<=4; end
			8065: begin bcd3<=8;bcd2<=0;bcd1<=6;bcd0<=5; end
			8066: begin bcd3<=8;bcd2<=0;bcd1<=6;bcd0<=6; end
			8067: begin bcd3<=8;bcd2<=0;bcd1<=6;bcd0<=7; end
			8068: begin bcd3<=8;bcd2<=0;bcd1<=6;bcd0<=8; end
			8069: begin bcd3<=8;bcd2<=0;bcd1<=6;bcd0<=9; end
			8070: begin bcd3<=8;bcd2<=0;bcd1<=7;bcd0<=0; end
			8071: begin bcd3<=8;bcd2<=0;bcd1<=7;bcd0<=1; end
			8072: begin bcd3<=8;bcd2<=0;bcd1<=7;bcd0<=2; end
			8073: begin bcd3<=8;bcd2<=0;bcd1<=7;bcd0<=3; end
			8074: begin bcd3<=8;bcd2<=0;bcd1<=7;bcd0<=4; end
			8075: begin bcd3<=8;bcd2<=0;bcd1<=7;bcd0<=5; end
			8076: begin bcd3<=8;bcd2<=0;bcd1<=7;bcd0<=6; end
			8077: begin bcd3<=8;bcd2<=0;bcd1<=7;bcd0<=7; end
			8078: begin bcd3<=8;bcd2<=0;bcd1<=7;bcd0<=8; end
			8079: begin bcd3<=8;bcd2<=0;bcd1<=7;bcd0<=9; end
			8080: begin bcd3<=8;bcd2<=0;bcd1<=8;bcd0<=0; end
			8081: begin bcd3<=8;bcd2<=0;bcd1<=8;bcd0<=1; end
			8082: begin bcd3<=8;bcd2<=0;bcd1<=8;bcd0<=2; end
			8083: begin bcd3<=8;bcd2<=0;bcd1<=8;bcd0<=3; end
			8084: begin bcd3<=8;bcd2<=0;bcd1<=8;bcd0<=4; end
			8085: begin bcd3<=8;bcd2<=0;bcd1<=8;bcd0<=5; end
			8086: begin bcd3<=8;bcd2<=0;bcd1<=8;bcd0<=6; end
			8087: begin bcd3<=8;bcd2<=0;bcd1<=8;bcd0<=7; end
			8088: begin bcd3<=8;bcd2<=0;bcd1<=8;bcd0<=8; end
			8089: begin bcd3<=8;bcd2<=0;bcd1<=8;bcd0<=9; end
			8090: begin bcd3<=8;bcd2<=0;bcd1<=9;bcd0<=0; end
			8091: begin bcd3<=8;bcd2<=0;bcd1<=9;bcd0<=1; end
			8092: begin bcd3<=8;bcd2<=0;bcd1<=9;bcd0<=2; end
			8093: begin bcd3<=8;bcd2<=0;bcd1<=9;bcd0<=3; end
			8094: begin bcd3<=8;bcd2<=0;bcd1<=9;bcd0<=4; end
			8095: begin bcd3<=8;bcd2<=0;bcd1<=9;bcd0<=5; end
			8096: begin bcd3<=8;bcd2<=0;bcd1<=9;bcd0<=6; end
			8097: begin bcd3<=8;bcd2<=0;bcd1<=9;bcd0<=7; end
			8098: begin bcd3<=8;bcd2<=0;bcd1<=9;bcd0<=8; end
			8099: begin bcd3<=8;bcd2<=0;bcd1<=9;bcd0<=9; end
			8100: begin bcd3<=8;bcd2<=1;bcd1<=0;bcd0<=0; end
			8101: begin bcd3<=8;bcd2<=1;bcd1<=0;bcd0<=1; end
			8102: begin bcd3<=8;bcd2<=1;bcd1<=0;bcd0<=2; end
			8103: begin bcd3<=8;bcd2<=1;bcd1<=0;bcd0<=3; end
			8104: begin bcd3<=8;bcd2<=1;bcd1<=0;bcd0<=4; end
			8105: begin bcd3<=8;bcd2<=1;bcd1<=0;bcd0<=5; end
			8106: begin bcd3<=8;bcd2<=1;bcd1<=0;bcd0<=6; end
			8107: begin bcd3<=8;bcd2<=1;bcd1<=0;bcd0<=7; end
			8108: begin bcd3<=8;bcd2<=1;bcd1<=0;bcd0<=8; end
			8109: begin bcd3<=8;bcd2<=1;bcd1<=0;bcd0<=9; end
			8110: begin bcd3<=8;bcd2<=1;bcd1<=1;bcd0<=0; end
			8111: begin bcd3<=8;bcd2<=1;bcd1<=1;bcd0<=1; end
			8112: begin bcd3<=8;bcd2<=1;bcd1<=1;bcd0<=2; end
			8113: begin bcd3<=8;bcd2<=1;bcd1<=1;bcd0<=3; end
			8114: begin bcd3<=8;bcd2<=1;bcd1<=1;bcd0<=4; end
			8115: begin bcd3<=8;bcd2<=1;bcd1<=1;bcd0<=5; end
			8116: begin bcd3<=8;bcd2<=1;bcd1<=1;bcd0<=6; end
			8117: begin bcd3<=8;bcd2<=1;bcd1<=1;bcd0<=7; end
			8118: begin bcd3<=8;bcd2<=1;bcd1<=1;bcd0<=8; end
			8119: begin bcd3<=8;bcd2<=1;bcd1<=1;bcd0<=9; end
			8120: begin bcd3<=8;bcd2<=1;bcd1<=2;bcd0<=0; end
			8121: begin bcd3<=8;bcd2<=1;bcd1<=2;bcd0<=1; end
			8122: begin bcd3<=8;bcd2<=1;bcd1<=2;bcd0<=2; end
			8123: begin bcd3<=8;bcd2<=1;bcd1<=2;bcd0<=3; end
			8124: begin bcd3<=8;bcd2<=1;bcd1<=2;bcd0<=4; end
			8125: begin bcd3<=8;bcd2<=1;bcd1<=2;bcd0<=5; end
			8126: begin bcd3<=8;bcd2<=1;bcd1<=2;bcd0<=6; end
			8127: begin bcd3<=8;bcd2<=1;bcd1<=2;bcd0<=7; end
			8128: begin bcd3<=8;bcd2<=1;bcd1<=2;bcd0<=8; end
			8129: begin bcd3<=8;bcd2<=1;bcd1<=2;bcd0<=9; end
			8130: begin bcd3<=8;bcd2<=1;bcd1<=3;bcd0<=0; end
			8131: begin bcd3<=8;bcd2<=1;bcd1<=3;bcd0<=1; end
			8132: begin bcd3<=8;bcd2<=1;bcd1<=3;bcd0<=2; end
			8133: begin bcd3<=8;bcd2<=1;bcd1<=3;bcd0<=3; end
			8134: begin bcd3<=8;bcd2<=1;bcd1<=3;bcd0<=4; end
			8135: begin bcd3<=8;bcd2<=1;bcd1<=3;bcd0<=5; end
			8136: begin bcd3<=8;bcd2<=1;bcd1<=3;bcd0<=6; end
			8137: begin bcd3<=8;bcd2<=1;bcd1<=3;bcd0<=7; end
			8138: begin bcd3<=8;bcd2<=1;bcd1<=3;bcd0<=8; end
			8139: begin bcd3<=8;bcd2<=1;bcd1<=3;bcd0<=9; end
			8140: begin bcd3<=8;bcd2<=1;bcd1<=4;bcd0<=0; end
			8141: begin bcd3<=8;bcd2<=1;bcd1<=4;bcd0<=1; end
			8142: begin bcd3<=8;bcd2<=1;bcd1<=4;bcd0<=2; end
			8143: begin bcd3<=8;bcd2<=1;bcd1<=4;bcd0<=3; end
			8144: begin bcd3<=8;bcd2<=1;bcd1<=4;bcd0<=4; end
			8145: begin bcd3<=8;bcd2<=1;bcd1<=4;bcd0<=5; end
			8146: begin bcd3<=8;bcd2<=1;bcd1<=4;bcd0<=6; end
			8147: begin bcd3<=8;bcd2<=1;bcd1<=4;bcd0<=7; end
			8148: begin bcd3<=8;bcd2<=1;bcd1<=4;bcd0<=8; end
			8149: begin bcd3<=8;bcd2<=1;bcd1<=4;bcd0<=9; end
			8150: begin bcd3<=8;bcd2<=1;bcd1<=5;bcd0<=0; end
			8151: begin bcd3<=8;bcd2<=1;bcd1<=5;bcd0<=1; end
			8152: begin bcd3<=8;bcd2<=1;bcd1<=5;bcd0<=2; end
			8153: begin bcd3<=8;bcd2<=1;bcd1<=5;bcd0<=3; end
			8154: begin bcd3<=8;bcd2<=1;bcd1<=5;bcd0<=4; end
			8155: begin bcd3<=8;bcd2<=1;bcd1<=5;bcd0<=5; end
			8156: begin bcd3<=8;bcd2<=1;bcd1<=5;bcd0<=6; end
			8157: begin bcd3<=8;bcd2<=1;bcd1<=5;bcd0<=7; end
			8158: begin bcd3<=8;bcd2<=1;bcd1<=5;bcd0<=8; end
			8159: begin bcd3<=8;bcd2<=1;bcd1<=5;bcd0<=9; end
			8160: begin bcd3<=8;bcd2<=1;bcd1<=6;bcd0<=0; end
			8161: begin bcd3<=8;bcd2<=1;bcd1<=6;bcd0<=1; end
			8162: begin bcd3<=8;bcd2<=1;bcd1<=6;bcd0<=2; end
			8163: begin bcd3<=8;bcd2<=1;bcd1<=6;bcd0<=3; end
			8164: begin bcd3<=8;bcd2<=1;bcd1<=6;bcd0<=4; end
			8165: begin bcd3<=8;bcd2<=1;bcd1<=6;bcd0<=5; end
			8166: begin bcd3<=8;bcd2<=1;bcd1<=6;bcd0<=6; end
			8167: begin bcd3<=8;bcd2<=1;bcd1<=6;bcd0<=7; end
			8168: begin bcd3<=8;bcd2<=1;bcd1<=6;bcd0<=8; end
			8169: begin bcd3<=8;bcd2<=1;bcd1<=6;bcd0<=9; end
			8170: begin bcd3<=8;bcd2<=1;bcd1<=7;bcd0<=0; end
			8171: begin bcd3<=8;bcd2<=1;bcd1<=7;bcd0<=1; end
			8172: begin bcd3<=8;bcd2<=1;bcd1<=7;bcd0<=2; end
			8173: begin bcd3<=8;bcd2<=1;bcd1<=7;bcd0<=3; end
			8174: begin bcd3<=8;bcd2<=1;bcd1<=7;bcd0<=4; end
			8175: begin bcd3<=8;bcd2<=1;bcd1<=7;bcd0<=5; end
			8176: begin bcd3<=8;bcd2<=1;bcd1<=7;bcd0<=6; end
			8177: begin bcd3<=8;bcd2<=1;bcd1<=7;bcd0<=7; end
			8178: begin bcd3<=8;bcd2<=1;bcd1<=7;bcd0<=8; end
			8179: begin bcd3<=8;bcd2<=1;bcd1<=7;bcd0<=9; end
			8180: begin bcd3<=8;bcd2<=1;bcd1<=8;bcd0<=0; end
			8181: begin bcd3<=8;bcd2<=1;bcd1<=8;bcd0<=1; end
			8182: begin bcd3<=8;bcd2<=1;bcd1<=8;bcd0<=2; end
			8183: begin bcd3<=8;bcd2<=1;bcd1<=8;bcd0<=3; end
			8184: begin bcd3<=8;bcd2<=1;bcd1<=8;bcd0<=4; end
			8185: begin bcd3<=8;bcd2<=1;bcd1<=8;bcd0<=5; end
			8186: begin bcd3<=8;bcd2<=1;bcd1<=8;bcd0<=6; end
			8187: begin bcd3<=8;bcd2<=1;bcd1<=8;bcd0<=7; end
			8188: begin bcd3<=8;bcd2<=1;bcd1<=8;bcd0<=8; end
			8189: begin bcd3<=8;bcd2<=1;bcd1<=8;bcd0<=9; end
			8190: begin bcd3<=8;bcd2<=1;bcd1<=9;bcd0<=0; end
			8191: begin bcd3<=8;bcd2<=1;bcd1<=9;bcd0<=1; end
			8192: begin bcd3<=8;bcd2<=1;bcd1<=9;bcd0<=2; end
			8193: begin bcd3<=8;bcd2<=1;bcd1<=9;bcd0<=3; end
			8194: begin bcd3<=8;bcd2<=1;bcd1<=9;bcd0<=4; end
			8195: begin bcd3<=8;bcd2<=1;bcd1<=9;bcd0<=5; end
			8196: begin bcd3<=8;bcd2<=1;bcd1<=9;bcd0<=6; end
			8197: begin bcd3<=8;bcd2<=1;bcd1<=9;bcd0<=7; end
			8198: begin bcd3<=8;bcd2<=1;bcd1<=9;bcd0<=8; end
			8199: begin bcd3<=8;bcd2<=1;bcd1<=9;bcd0<=9; end
			8200: begin bcd3<=8;bcd2<=2;bcd1<=0;bcd0<=0; end
			8201: begin bcd3<=8;bcd2<=2;bcd1<=0;bcd0<=1; end
			8202: begin bcd3<=8;bcd2<=2;bcd1<=0;bcd0<=2; end
			8203: begin bcd3<=8;bcd2<=2;bcd1<=0;bcd0<=3; end
			8204: begin bcd3<=8;bcd2<=2;bcd1<=0;bcd0<=4; end
			8205: begin bcd3<=8;bcd2<=2;bcd1<=0;bcd0<=5; end
			8206: begin bcd3<=8;bcd2<=2;bcd1<=0;bcd0<=6; end
			8207: begin bcd3<=8;bcd2<=2;bcd1<=0;bcd0<=7; end
			8208: begin bcd3<=8;bcd2<=2;bcd1<=0;bcd0<=8; end
			8209: begin bcd3<=8;bcd2<=2;bcd1<=0;bcd0<=9; end
			8210: begin bcd3<=8;bcd2<=2;bcd1<=1;bcd0<=0; end
			8211: begin bcd3<=8;bcd2<=2;bcd1<=1;bcd0<=1; end
			8212: begin bcd3<=8;bcd2<=2;bcd1<=1;bcd0<=2; end
			8213: begin bcd3<=8;bcd2<=2;bcd1<=1;bcd0<=3; end
			8214: begin bcd3<=8;bcd2<=2;bcd1<=1;bcd0<=4; end
			8215: begin bcd3<=8;bcd2<=2;bcd1<=1;bcd0<=5; end
			8216: begin bcd3<=8;bcd2<=2;bcd1<=1;bcd0<=6; end
			8217: begin bcd3<=8;bcd2<=2;bcd1<=1;bcd0<=7; end
			8218: begin bcd3<=8;bcd2<=2;bcd1<=1;bcd0<=8; end
			8219: begin bcd3<=8;bcd2<=2;bcd1<=1;bcd0<=9; end
			8220: begin bcd3<=8;bcd2<=2;bcd1<=2;bcd0<=0; end
			8221: begin bcd3<=8;bcd2<=2;bcd1<=2;bcd0<=1; end
			8222: begin bcd3<=8;bcd2<=2;bcd1<=2;bcd0<=2; end
			8223: begin bcd3<=8;bcd2<=2;bcd1<=2;bcd0<=3; end
			8224: begin bcd3<=8;bcd2<=2;bcd1<=2;bcd0<=4; end
			8225: begin bcd3<=8;bcd2<=2;bcd1<=2;bcd0<=5; end
			8226: begin bcd3<=8;bcd2<=2;bcd1<=2;bcd0<=6; end
			8227: begin bcd3<=8;bcd2<=2;bcd1<=2;bcd0<=7; end
			8228: begin bcd3<=8;bcd2<=2;bcd1<=2;bcd0<=8; end
			8229: begin bcd3<=8;bcd2<=2;bcd1<=2;bcd0<=9; end
			8230: begin bcd3<=8;bcd2<=2;bcd1<=3;bcd0<=0; end
			8231: begin bcd3<=8;bcd2<=2;bcd1<=3;bcd0<=1; end
			8232: begin bcd3<=8;bcd2<=2;bcd1<=3;bcd0<=2; end
			8233: begin bcd3<=8;bcd2<=2;bcd1<=3;bcd0<=3; end
			8234: begin bcd3<=8;bcd2<=2;bcd1<=3;bcd0<=4; end
			8235: begin bcd3<=8;bcd2<=2;bcd1<=3;bcd0<=5; end
			8236: begin bcd3<=8;bcd2<=2;bcd1<=3;bcd0<=6; end
			8237: begin bcd3<=8;bcd2<=2;bcd1<=3;bcd0<=7; end
			8238: begin bcd3<=8;bcd2<=2;bcd1<=3;bcd0<=8; end
			8239: begin bcd3<=8;bcd2<=2;bcd1<=3;bcd0<=9; end
			8240: begin bcd3<=8;bcd2<=2;bcd1<=4;bcd0<=0; end
			8241: begin bcd3<=8;bcd2<=2;bcd1<=4;bcd0<=1; end
			8242: begin bcd3<=8;bcd2<=2;bcd1<=4;bcd0<=2; end
			8243: begin bcd3<=8;bcd2<=2;bcd1<=4;bcd0<=3; end
			8244: begin bcd3<=8;bcd2<=2;bcd1<=4;bcd0<=4; end
			8245: begin bcd3<=8;bcd2<=2;bcd1<=4;bcd0<=5; end
			8246: begin bcd3<=8;bcd2<=2;bcd1<=4;bcd0<=6; end
			8247: begin bcd3<=8;bcd2<=2;bcd1<=4;bcd0<=7; end
			8248: begin bcd3<=8;bcd2<=2;bcd1<=4;bcd0<=8; end
			8249: begin bcd3<=8;bcd2<=2;bcd1<=4;bcd0<=9; end
			8250: begin bcd3<=8;bcd2<=2;bcd1<=5;bcd0<=0; end
			8251: begin bcd3<=8;bcd2<=2;bcd1<=5;bcd0<=1; end
			8252: begin bcd3<=8;bcd2<=2;bcd1<=5;bcd0<=2; end
			8253: begin bcd3<=8;bcd2<=2;bcd1<=5;bcd0<=3; end
			8254: begin bcd3<=8;bcd2<=2;bcd1<=5;bcd0<=4; end
			8255: begin bcd3<=8;bcd2<=2;bcd1<=5;bcd0<=5; end
			8256: begin bcd3<=8;bcd2<=2;bcd1<=5;bcd0<=6; end
			8257: begin bcd3<=8;bcd2<=2;bcd1<=5;bcd0<=7; end
			8258: begin bcd3<=8;bcd2<=2;bcd1<=5;bcd0<=8; end
			8259: begin bcd3<=8;bcd2<=2;bcd1<=5;bcd0<=9; end
			8260: begin bcd3<=8;bcd2<=2;bcd1<=6;bcd0<=0; end
			8261: begin bcd3<=8;bcd2<=2;bcd1<=6;bcd0<=1; end
			8262: begin bcd3<=8;bcd2<=2;bcd1<=6;bcd0<=2; end
			8263: begin bcd3<=8;bcd2<=2;bcd1<=6;bcd0<=3; end
			8264: begin bcd3<=8;bcd2<=2;bcd1<=6;bcd0<=4; end
			8265: begin bcd3<=8;bcd2<=2;bcd1<=6;bcd0<=5; end
			8266: begin bcd3<=8;bcd2<=2;bcd1<=6;bcd0<=6; end
			8267: begin bcd3<=8;bcd2<=2;bcd1<=6;bcd0<=7; end
			8268: begin bcd3<=8;bcd2<=2;bcd1<=6;bcd0<=8; end
			8269: begin bcd3<=8;bcd2<=2;bcd1<=6;bcd0<=9; end
			8270: begin bcd3<=8;bcd2<=2;bcd1<=7;bcd0<=0; end
			8271: begin bcd3<=8;bcd2<=2;bcd1<=7;bcd0<=1; end
			8272: begin bcd3<=8;bcd2<=2;bcd1<=7;bcd0<=2; end
			8273: begin bcd3<=8;bcd2<=2;bcd1<=7;bcd0<=3; end
			8274: begin bcd3<=8;bcd2<=2;bcd1<=7;bcd0<=4; end
			8275: begin bcd3<=8;bcd2<=2;bcd1<=7;bcd0<=5; end
			8276: begin bcd3<=8;bcd2<=2;bcd1<=7;bcd0<=6; end
			8277: begin bcd3<=8;bcd2<=2;bcd1<=7;bcd0<=7; end
			8278: begin bcd3<=8;bcd2<=2;bcd1<=7;bcd0<=8; end
			8279: begin bcd3<=8;bcd2<=2;bcd1<=7;bcd0<=9; end
			8280: begin bcd3<=8;bcd2<=2;bcd1<=8;bcd0<=0; end
			8281: begin bcd3<=8;bcd2<=2;bcd1<=8;bcd0<=1; end
			8282: begin bcd3<=8;bcd2<=2;bcd1<=8;bcd0<=2; end
			8283: begin bcd3<=8;bcd2<=2;bcd1<=8;bcd0<=3; end
			8284: begin bcd3<=8;bcd2<=2;bcd1<=8;bcd0<=4; end
			8285: begin bcd3<=8;bcd2<=2;bcd1<=8;bcd0<=5; end
			8286: begin bcd3<=8;bcd2<=2;bcd1<=8;bcd0<=6; end
			8287: begin bcd3<=8;bcd2<=2;bcd1<=8;bcd0<=7; end
			8288: begin bcd3<=8;bcd2<=2;bcd1<=8;bcd0<=8; end
			8289: begin bcd3<=8;bcd2<=2;bcd1<=8;bcd0<=9; end
			8290: begin bcd3<=8;bcd2<=2;bcd1<=9;bcd0<=0; end
			8291: begin bcd3<=8;bcd2<=2;bcd1<=9;bcd0<=1; end
			8292: begin bcd3<=8;bcd2<=2;bcd1<=9;bcd0<=2; end
			8293: begin bcd3<=8;bcd2<=2;bcd1<=9;bcd0<=3; end
			8294: begin bcd3<=8;bcd2<=2;bcd1<=9;bcd0<=4; end
			8295: begin bcd3<=8;bcd2<=2;bcd1<=9;bcd0<=5; end
			8296: begin bcd3<=8;bcd2<=2;bcd1<=9;bcd0<=6; end
			8297: begin bcd3<=8;bcd2<=2;bcd1<=9;bcd0<=7; end
			8298: begin bcd3<=8;bcd2<=2;bcd1<=9;bcd0<=8; end
			8299: begin bcd3<=8;bcd2<=2;bcd1<=9;bcd0<=9; end
			8300: begin bcd3<=8;bcd2<=3;bcd1<=0;bcd0<=0; end
			8301: begin bcd3<=8;bcd2<=3;bcd1<=0;bcd0<=1; end
			8302: begin bcd3<=8;bcd2<=3;bcd1<=0;bcd0<=2; end
			8303: begin bcd3<=8;bcd2<=3;bcd1<=0;bcd0<=3; end
			8304: begin bcd3<=8;bcd2<=3;bcd1<=0;bcd0<=4; end
			8305: begin bcd3<=8;bcd2<=3;bcd1<=0;bcd0<=5; end
			8306: begin bcd3<=8;bcd2<=3;bcd1<=0;bcd0<=6; end
			8307: begin bcd3<=8;bcd2<=3;bcd1<=0;bcd0<=7; end
			8308: begin bcd3<=8;bcd2<=3;bcd1<=0;bcd0<=8; end
			8309: begin bcd3<=8;bcd2<=3;bcd1<=0;bcd0<=9; end
			8310: begin bcd3<=8;bcd2<=3;bcd1<=1;bcd0<=0; end
			8311: begin bcd3<=8;bcd2<=3;bcd1<=1;bcd0<=1; end
			8312: begin bcd3<=8;bcd2<=3;bcd1<=1;bcd0<=2; end
			8313: begin bcd3<=8;bcd2<=3;bcd1<=1;bcd0<=3; end
			8314: begin bcd3<=8;bcd2<=3;bcd1<=1;bcd0<=4; end
			8315: begin bcd3<=8;bcd2<=3;bcd1<=1;bcd0<=5; end
			8316: begin bcd3<=8;bcd2<=3;bcd1<=1;bcd0<=6; end
			8317: begin bcd3<=8;bcd2<=3;bcd1<=1;bcd0<=7; end
			8318: begin bcd3<=8;bcd2<=3;bcd1<=1;bcd0<=8; end
			8319: begin bcd3<=8;bcd2<=3;bcd1<=1;bcd0<=9; end
			8320: begin bcd3<=8;bcd2<=3;bcd1<=2;bcd0<=0; end
			8321: begin bcd3<=8;bcd2<=3;bcd1<=2;bcd0<=1; end
			8322: begin bcd3<=8;bcd2<=3;bcd1<=2;bcd0<=2; end
			8323: begin bcd3<=8;bcd2<=3;bcd1<=2;bcd0<=3; end
			8324: begin bcd3<=8;bcd2<=3;bcd1<=2;bcd0<=4; end
			8325: begin bcd3<=8;bcd2<=3;bcd1<=2;bcd0<=5; end
			8326: begin bcd3<=8;bcd2<=3;bcd1<=2;bcd0<=6; end
			8327: begin bcd3<=8;bcd2<=3;bcd1<=2;bcd0<=7; end
			8328: begin bcd3<=8;bcd2<=3;bcd1<=2;bcd0<=8; end
			8329: begin bcd3<=8;bcd2<=3;bcd1<=2;bcd0<=9; end
			8330: begin bcd3<=8;bcd2<=3;bcd1<=3;bcd0<=0; end
			8331: begin bcd3<=8;bcd2<=3;bcd1<=3;bcd0<=1; end
			8332: begin bcd3<=8;bcd2<=3;bcd1<=3;bcd0<=2; end
			8333: begin bcd3<=8;bcd2<=3;bcd1<=3;bcd0<=3; end
			8334: begin bcd3<=8;bcd2<=3;bcd1<=3;bcd0<=4; end
			8335: begin bcd3<=8;bcd2<=3;bcd1<=3;bcd0<=5; end
			8336: begin bcd3<=8;bcd2<=3;bcd1<=3;bcd0<=6; end
			8337: begin bcd3<=8;bcd2<=3;bcd1<=3;bcd0<=7; end
			8338: begin bcd3<=8;bcd2<=3;bcd1<=3;bcd0<=8; end
			8339: begin bcd3<=8;bcd2<=3;bcd1<=3;bcd0<=9; end
			8340: begin bcd3<=8;bcd2<=3;bcd1<=4;bcd0<=0; end
			8341: begin bcd3<=8;bcd2<=3;bcd1<=4;bcd0<=1; end
			8342: begin bcd3<=8;bcd2<=3;bcd1<=4;bcd0<=2; end
			8343: begin bcd3<=8;bcd2<=3;bcd1<=4;bcd0<=3; end
			8344: begin bcd3<=8;bcd2<=3;bcd1<=4;bcd0<=4; end
			8345: begin bcd3<=8;bcd2<=3;bcd1<=4;bcd0<=5; end
			8346: begin bcd3<=8;bcd2<=3;bcd1<=4;bcd0<=6; end
			8347: begin bcd3<=8;bcd2<=3;bcd1<=4;bcd0<=7; end
			8348: begin bcd3<=8;bcd2<=3;bcd1<=4;bcd0<=8; end
			8349: begin bcd3<=8;bcd2<=3;bcd1<=4;bcd0<=9; end
			8350: begin bcd3<=8;bcd2<=3;bcd1<=5;bcd0<=0; end
			8351: begin bcd3<=8;bcd2<=3;bcd1<=5;bcd0<=1; end
			8352: begin bcd3<=8;bcd2<=3;bcd1<=5;bcd0<=2; end
			8353: begin bcd3<=8;bcd2<=3;bcd1<=5;bcd0<=3; end
			8354: begin bcd3<=8;bcd2<=3;bcd1<=5;bcd0<=4; end
			8355: begin bcd3<=8;bcd2<=3;bcd1<=5;bcd0<=5; end
			8356: begin bcd3<=8;bcd2<=3;bcd1<=5;bcd0<=6; end
			8357: begin bcd3<=8;bcd2<=3;bcd1<=5;bcd0<=7; end
			8358: begin bcd3<=8;bcd2<=3;bcd1<=5;bcd0<=8; end
			8359: begin bcd3<=8;bcd2<=3;bcd1<=5;bcd0<=9; end
			8360: begin bcd3<=8;bcd2<=3;bcd1<=6;bcd0<=0; end
			8361: begin bcd3<=8;bcd2<=3;bcd1<=6;bcd0<=1; end
			8362: begin bcd3<=8;bcd2<=3;bcd1<=6;bcd0<=2; end
			8363: begin bcd3<=8;bcd2<=3;bcd1<=6;bcd0<=3; end
			8364: begin bcd3<=8;bcd2<=3;bcd1<=6;bcd0<=4; end
			8365: begin bcd3<=8;bcd2<=3;bcd1<=6;bcd0<=5; end
			8366: begin bcd3<=8;bcd2<=3;bcd1<=6;bcd0<=6; end
			8367: begin bcd3<=8;bcd2<=3;bcd1<=6;bcd0<=7; end
			8368: begin bcd3<=8;bcd2<=3;bcd1<=6;bcd0<=8; end
			8369: begin bcd3<=8;bcd2<=3;bcd1<=6;bcd0<=9; end
			8370: begin bcd3<=8;bcd2<=3;bcd1<=7;bcd0<=0; end
			8371: begin bcd3<=8;bcd2<=3;bcd1<=7;bcd0<=1; end
			8372: begin bcd3<=8;bcd2<=3;bcd1<=7;bcd0<=2; end
			8373: begin bcd3<=8;bcd2<=3;bcd1<=7;bcd0<=3; end
			8374: begin bcd3<=8;bcd2<=3;bcd1<=7;bcd0<=4; end
			8375: begin bcd3<=8;bcd2<=3;bcd1<=7;bcd0<=5; end
			8376: begin bcd3<=8;bcd2<=3;bcd1<=7;bcd0<=6; end
			8377: begin bcd3<=8;bcd2<=3;bcd1<=7;bcd0<=7; end
			8378: begin bcd3<=8;bcd2<=3;bcd1<=7;bcd0<=8; end
			8379: begin bcd3<=8;bcd2<=3;bcd1<=7;bcd0<=9; end
			8380: begin bcd3<=8;bcd2<=3;bcd1<=8;bcd0<=0; end
			8381: begin bcd3<=8;bcd2<=3;bcd1<=8;bcd0<=1; end
			8382: begin bcd3<=8;bcd2<=3;bcd1<=8;bcd0<=2; end
			8383: begin bcd3<=8;bcd2<=3;bcd1<=8;bcd0<=3; end
			8384: begin bcd3<=8;bcd2<=3;bcd1<=8;bcd0<=4; end
			8385: begin bcd3<=8;bcd2<=3;bcd1<=8;bcd0<=5; end
			8386: begin bcd3<=8;bcd2<=3;bcd1<=8;bcd0<=6; end
			8387: begin bcd3<=8;bcd2<=3;bcd1<=8;bcd0<=7; end
			8388: begin bcd3<=8;bcd2<=3;bcd1<=8;bcd0<=8; end
			8389: begin bcd3<=8;bcd2<=3;bcd1<=8;bcd0<=9; end
			8390: begin bcd3<=8;bcd2<=3;bcd1<=9;bcd0<=0; end
			8391: begin bcd3<=8;bcd2<=3;bcd1<=9;bcd0<=1; end
			8392: begin bcd3<=8;bcd2<=3;bcd1<=9;bcd0<=2; end
			8393: begin bcd3<=8;bcd2<=3;bcd1<=9;bcd0<=3; end
			8394: begin bcd3<=8;bcd2<=3;bcd1<=9;bcd0<=4; end
			8395: begin bcd3<=8;bcd2<=3;bcd1<=9;bcd0<=5; end
			8396: begin bcd3<=8;bcd2<=3;bcd1<=9;bcd0<=6; end
			8397: begin bcd3<=8;bcd2<=3;bcd1<=9;bcd0<=7; end
			8398: begin bcd3<=8;bcd2<=3;bcd1<=9;bcd0<=8; end
			8399: begin bcd3<=8;bcd2<=3;bcd1<=9;bcd0<=9; end
			8400: begin bcd3<=8;bcd2<=4;bcd1<=0;bcd0<=0; end
			8401: begin bcd3<=8;bcd2<=4;bcd1<=0;bcd0<=1; end
			8402: begin bcd3<=8;bcd2<=4;bcd1<=0;bcd0<=2; end
			8403: begin bcd3<=8;bcd2<=4;bcd1<=0;bcd0<=3; end
			8404: begin bcd3<=8;bcd2<=4;bcd1<=0;bcd0<=4; end
			8405: begin bcd3<=8;bcd2<=4;bcd1<=0;bcd0<=5; end
			8406: begin bcd3<=8;bcd2<=4;bcd1<=0;bcd0<=6; end
			8407: begin bcd3<=8;bcd2<=4;bcd1<=0;bcd0<=7; end
			8408: begin bcd3<=8;bcd2<=4;bcd1<=0;bcd0<=8; end
			8409: begin bcd3<=8;bcd2<=4;bcd1<=0;bcd0<=9; end
			8410: begin bcd3<=8;bcd2<=4;bcd1<=1;bcd0<=0; end
			8411: begin bcd3<=8;bcd2<=4;bcd1<=1;bcd0<=1; end
			8412: begin bcd3<=8;bcd2<=4;bcd1<=1;bcd0<=2; end
			8413: begin bcd3<=8;bcd2<=4;bcd1<=1;bcd0<=3; end
			8414: begin bcd3<=8;bcd2<=4;bcd1<=1;bcd0<=4; end
			8415: begin bcd3<=8;bcd2<=4;bcd1<=1;bcd0<=5; end
			8416: begin bcd3<=8;bcd2<=4;bcd1<=1;bcd0<=6; end
			8417: begin bcd3<=8;bcd2<=4;bcd1<=1;bcd0<=7; end
			8418: begin bcd3<=8;bcd2<=4;bcd1<=1;bcd0<=8; end
			8419: begin bcd3<=8;bcd2<=4;bcd1<=1;bcd0<=9; end
			8420: begin bcd3<=8;bcd2<=4;bcd1<=2;bcd0<=0; end
			8421: begin bcd3<=8;bcd2<=4;bcd1<=2;bcd0<=1; end
			8422: begin bcd3<=8;bcd2<=4;bcd1<=2;bcd0<=2; end
			8423: begin bcd3<=8;bcd2<=4;bcd1<=2;bcd0<=3; end
			8424: begin bcd3<=8;bcd2<=4;bcd1<=2;bcd0<=4; end
			8425: begin bcd3<=8;bcd2<=4;bcd1<=2;bcd0<=5; end
			8426: begin bcd3<=8;bcd2<=4;bcd1<=2;bcd0<=6; end
			8427: begin bcd3<=8;bcd2<=4;bcd1<=2;bcd0<=7; end
			8428: begin bcd3<=8;bcd2<=4;bcd1<=2;bcd0<=8; end
			8429: begin bcd3<=8;bcd2<=4;bcd1<=2;bcd0<=9; end
			8430: begin bcd3<=8;bcd2<=4;bcd1<=3;bcd0<=0; end
			8431: begin bcd3<=8;bcd2<=4;bcd1<=3;bcd0<=1; end
			8432: begin bcd3<=8;bcd2<=4;bcd1<=3;bcd0<=2; end
			8433: begin bcd3<=8;bcd2<=4;bcd1<=3;bcd0<=3; end
			8434: begin bcd3<=8;bcd2<=4;bcd1<=3;bcd0<=4; end
			8435: begin bcd3<=8;bcd2<=4;bcd1<=3;bcd0<=5; end
			8436: begin bcd3<=8;bcd2<=4;bcd1<=3;bcd0<=6; end
			8437: begin bcd3<=8;bcd2<=4;bcd1<=3;bcd0<=7; end
			8438: begin bcd3<=8;bcd2<=4;bcd1<=3;bcd0<=8; end
			8439: begin bcd3<=8;bcd2<=4;bcd1<=3;bcd0<=9; end
			8440: begin bcd3<=8;bcd2<=4;bcd1<=4;bcd0<=0; end
			8441: begin bcd3<=8;bcd2<=4;bcd1<=4;bcd0<=1; end
			8442: begin bcd3<=8;bcd2<=4;bcd1<=4;bcd0<=2; end
			8443: begin bcd3<=8;bcd2<=4;bcd1<=4;bcd0<=3; end
			8444: begin bcd3<=8;bcd2<=4;bcd1<=4;bcd0<=4; end
			8445: begin bcd3<=8;bcd2<=4;bcd1<=4;bcd0<=5; end
			8446: begin bcd3<=8;bcd2<=4;bcd1<=4;bcd0<=6; end
			8447: begin bcd3<=8;bcd2<=4;bcd1<=4;bcd0<=7; end
			8448: begin bcd3<=8;bcd2<=4;bcd1<=4;bcd0<=8; end
			8449: begin bcd3<=8;bcd2<=4;bcd1<=4;bcd0<=9; end
			8450: begin bcd3<=8;bcd2<=4;bcd1<=5;bcd0<=0; end
			8451: begin bcd3<=8;bcd2<=4;bcd1<=5;bcd0<=1; end
			8452: begin bcd3<=8;bcd2<=4;bcd1<=5;bcd0<=2; end
			8453: begin bcd3<=8;bcd2<=4;bcd1<=5;bcd0<=3; end
			8454: begin bcd3<=8;bcd2<=4;bcd1<=5;bcd0<=4; end
			8455: begin bcd3<=8;bcd2<=4;bcd1<=5;bcd0<=5; end
			8456: begin bcd3<=8;bcd2<=4;bcd1<=5;bcd0<=6; end
			8457: begin bcd3<=8;bcd2<=4;bcd1<=5;bcd0<=7; end
			8458: begin bcd3<=8;bcd2<=4;bcd1<=5;bcd0<=8; end
			8459: begin bcd3<=8;bcd2<=4;bcd1<=5;bcd0<=9; end
			8460: begin bcd3<=8;bcd2<=4;bcd1<=6;bcd0<=0; end
			8461: begin bcd3<=8;bcd2<=4;bcd1<=6;bcd0<=1; end
			8462: begin bcd3<=8;bcd2<=4;bcd1<=6;bcd0<=2; end
			8463: begin bcd3<=8;bcd2<=4;bcd1<=6;bcd0<=3; end
			8464: begin bcd3<=8;bcd2<=4;bcd1<=6;bcd0<=4; end
			8465: begin bcd3<=8;bcd2<=4;bcd1<=6;bcd0<=5; end
			8466: begin bcd3<=8;bcd2<=4;bcd1<=6;bcd0<=6; end
			8467: begin bcd3<=8;bcd2<=4;bcd1<=6;bcd0<=7; end
			8468: begin bcd3<=8;bcd2<=4;bcd1<=6;bcd0<=8; end
			8469: begin bcd3<=8;bcd2<=4;bcd1<=6;bcd0<=9; end
			8470: begin bcd3<=8;bcd2<=4;bcd1<=7;bcd0<=0; end
			8471: begin bcd3<=8;bcd2<=4;bcd1<=7;bcd0<=1; end
			8472: begin bcd3<=8;bcd2<=4;bcd1<=7;bcd0<=2; end
			8473: begin bcd3<=8;bcd2<=4;bcd1<=7;bcd0<=3; end
			8474: begin bcd3<=8;bcd2<=4;bcd1<=7;bcd0<=4; end
			8475: begin bcd3<=8;bcd2<=4;bcd1<=7;bcd0<=5; end
			8476: begin bcd3<=8;bcd2<=4;bcd1<=7;bcd0<=6; end
			8477: begin bcd3<=8;bcd2<=4;bcd1<=7;bcd0<=7; end
			8478: begin bcd3<=8;bcd2<=4;bcd1<=7;bcd0<=8; end
			8479: begin bcd3<=8;bcd2<=4;bcd1<=7;bcd0<=9; end
			8480: begin bcd3<=8;bcd2<=4;bcd1<=8;bcd0<=0; end
			8481: begin bcd3<=8;bcd2<=4;bcd1<=8;bcd0<=1; end
			8482: begin bcd3<=8;bcd2<=4;bcd1<=8;bcd0<=2; end
			8483: begin bcd3<=8;bcd2<=4;bcd1<=8;bcd0<=3; end
			8484: begin bcd3<=8;bcd2<=4;bcd1<=8;bcd0<=4; end
			8485: begin bcd3<=8;bcd2<=4;bcd1<=8;bcd0<=5; end
			8486: begin bcd3<=8;bcd2<=4;bcd1<=8;bcd0<=6; end
			8487: begin bcd3<=8;bcd2<=4;bcd1<=8;bcd0<=7; end
			8488: begin bcd3<=8;bcd2<=4;bcd1<=8;bcd0<=8; end
			8489: begin bcd3<=8;bcd2<=4;bcd1<=8;bcd0<=9; end
			8490: begin bcd3<=8;bcd2<=4;bcd1<=9;bcd0<=0; end
			8491: begin bcd3<=8;bcd2<=4;bcd1<=9;bcd0<=1; end
			8492: begin bcd3<=8;bcd2<=4;bcd1<=9;bcd0<=2; end
			8493: begin bcd3<=8;bcd2<=4;bcd1<=9;bcd0<=3; end
			8494: begin bcd3<=8;bcd2<=4;bcd1<=9;bcd0<=4; end
			8495: begin bcd3<=8;bcd2<=4;bcd1<=9;bcd0<=5; end
			8496: begin bcd3<=8;bcd2<=4;bcd1<=9;bcd0<=6; end
			8497: begin bcd3<=8;bcd2<=4;bcd1<=9;bcd0<=7; end
			8498: begin bcd3<=8;bcd2<=4;bcd1<=9;bcd0<=8; end
			8499: begin bcd3<=8;bcd2<=4;bcd1<=9;bcd0<=9; end
			8500: begin bcd3<=8;bcd2<=5;bcd1<=0;bcd0<=0; end
			8501: begin bcd3<=8;bcd2<=5;bcd1<=0;bcd0<=1; end
			8502: begin bcd3<=8;bcd2<=5;bcd1<=0;bcd0<=2; end
			8503: begin bcd3<=8;bcd2<=5;bcd1<=0;bcd0<=3; end
			8504: begin bcd3<=8;bcd2<=5;bcd1<=0;bcd0<=4; end
			8505: begin bcd3<=8;bcd2<=5;bcd1<=0;bcd0<=5; end
			8506: begin bcd3<=8;bcd2<=5;bcd1<=0;bcd0<=6; end
			8507: begin bcd3<=8;bcd2<=5;bcd1<=0;bcd0<=7; end
			8508: begin bcd3<=8;bcd2<=5;bcd1<=0;bcd0<=8; end
			8509: begin bcd3<=8;bcd2<=5;bcd1<=0;bcd0<=9; end
			8510: begin bcd3<=8;bcd2<=5;bcd1<=1;bcd0<=0; end
			8511: begin bcd3<=8;bcd2<=5;bcd1<=1;bcd0<=1; end
			8512: begin bcd3<=8;bcd2<=5;bcd1<=1;bcd0<=2; end
			8513: begin bcd3<=8;bcd2<=5;bcd1<=1;bcd0<=3; end
			8514: begin bcd3<=8;bcd2<=5;bcd1<=1;bcd0<=4; end
			8515: begin bcd3<=8;bcd2<=5;bcd1<=1;bcd0<=5; end
			8516: begin bcd3<=8;bcd2<=5;bcd1<=1;bcd0<=6; end
			8517: begin bcd3<=8;bcd2<=5;bcd1<=1;bcd0<=7; end
			8518: begin bcd3<=8;bcd2<=5;bcd1<=1;bcd0<=8; end
			8519: begin bcd3<=8;bcd2<=5;bcd1<=1;bcd0<=9; end
			8520: begin bcd3<=8;bcd2<=5;bcd1<=2;bcd0<=0; end
			8521: begin bcd3<=8;bcd2<=5;bcd1<=2;bcd0<=1; end
			8522: begin bcd3<=8;bcd2<=5;bcd1<=2;bcd0<=2; end
			8523: begin bcd3<=8;bcd2<=5;bcd1<=2;bcd0<=3; end
			8524: begin bcd3<=8;bcd2<=5;bcd1<=2;bcd0<=4; end
			8525: begin bcd3<=8;bcd2<=5;bcd1<=2;bcd0<=5; end
			8526: begin bcd3<=8;bcd2<=5;bcd1<=2;bcd0<=6; end
			8527: begin bcd3<=8;bcd2<=5;bcd1<=2;bcd0<=7; end
			8528: begin bcd3<=8;bcd2<=5;bcd1<=2;bcd0<=8; end
			8529: begin bcd3<=8;bcd2<=5;bcd1<=2;bcd0<=9; end
			8530: begin bcd3<=8;bcd2<=5;bcd1<=3;bcd0<=0; end
			8531: begin bcd3<=8;bcd2<=5;bcd1<=3;bcd0<=1; end
			8532: begin bcd3<=8;bcd2<=5;bcd1<=3;bcd0<=2; end
			8533: begin bcd3<=8;bcd2<=5;bcd1<=3;bcd0<=3; end
			8534: begin bcd3<=8;bcd2<=5;bcd1<=3;bcd0<=4; end
			8535: begin bcd3<=8;bcd2<=5;bcd1<=3;bcd0<=5; end
			8536: begin bcd3<=8;bcd2<=5;bcd1<=3;bcd0<=6; end
			8537: begin bcd3<=8;bcd2<=5;bcd1<=3;bcd0<=7; end
			8538: begin bcd3<=8;bcd2<=5;bcd1<=3;bcd0<=8; end
			8539: begin bcd3<=8;bcd2<=5;bcd1<=3;bcd0<=9; end
			8540: begin bcd3<=8;bcd2<=5;bcd1<=4;bcd0<=0; end
			8541: begin bcd3<=8;bcd2<=5;bcd1<=4;bcd0<=1; end
			8542: begin bcd3<=8;bcd2<=5;bcd1<=4;bcd0<=2; end
			8543: begin bcd3<=8;bcd2<=5;bcd1<=4;bcd0<=3; end
			8544: begin bcd3<=8;bcd2<=5;bcd1<=4;bcd0<=4; end
			8545: begin bcd3<=8;bcd2<=5;bcd1<=4;bcd0<=5; end
			8546: begin bcd3<=8;bcd2<=5;bcd1<=4;bcd0<=6; end
			8547: begin bcd3<=8;bcd2<=5;bcd1<=4;bcd0<=7; end
			8548: begin bcd3<=8;bcd2<=5;bcd1<=4;bcd0<=8; end
			8549: begin bcd3<=8;bcd2<=5;bcd1<=4;bcd0<=9; end
			8550: begin bcd3<=8;bcd2<=5;bcd1<=5;bcd0<=0; end
			8551: begin bcd3<=8;bcd2<=5;bcd1<=5;bcd0<=1; end
			8552: begin bcd3<=8;bcd2<=5;bcd1<=5;bcd0<=2; end
			8553: begin bcd3<=8;bcd2<=5;bcd1<=5;bcd0<=3; end
			8554: begin bcd3<=8;bcd2<=5;bcd1<=5;bcd0<=4; end
			8555: begin bcd3<=8;bcd2<=5;bcd1<=5;bcd0<=5; end
			8556: begin bcd3<=8;bcd2<=5;bcd1<=5;bcd0<=6; end
			8557: begin bcd3<=8;bcd2<=5;bcd1<=5;bcd0<=7; end
			8558: begin bcd3<=8;bcd2<=5;bcd1<=5;bcd0<=8; end
			8559: begin bcd3<=8;bcd2<=5;bcd1<=5;bcd0<=9; end
			8560: begin bcd3<=8;bcd2<=5;bcd1<=6;bcd0<=0; end
			8561: begin bcd3<=8;bcd2<=5;bcd1<=6;bcd0<=1; end
			8562: begin bcd3<=8;bcd2<=5;bcd1<=6;bcd0<=2; end
			8563: begin bcd3<=8;bcd2<=5;bcd1<=6;bcd0<=3; end
			8564: begin bcd3<=8;bcd2<=5;bcd1<=6;bcd0<=4; end
			8565: begin bcd3<=8;bcd2<=5;bcd1<=6;bcd0<=5; end
			8566: begin bcd3<=8;bcd2<=5;bcd1<=6;bcd0<=6; end
			8567: begin bcd3<=8;bcd2<=5;bcd1<=6;bcd0<=7; end
			8568: begin bcd3<=8;bcd2<=5;bcd1<=6;bcd0<=8; end
			8569: begin bcd3<=8;bcd2<=5;bcd1<=6;bcd0<=9; end
			8570: begin bcd3<=8;bcd2<=5;bcd1<=7;bcd0<=0; end
			8571: begin bcd3<=8;bcd2<=5;bcd1<=7;bcd0<=1; end
			8572: begin bcd3<=8;bcd2<=5;bcd1<=7;bcd0<=2; end
			8573: begin bcd3<=8;bcd2<=5;bcd1<=7;bcd0<=3; end
			8574: begin bcd3<=8;bcd2<=5;bcd1<=7;bcd0<=4; end
			8575: begin bcd3<=8;bcd2<=5;bcd1<=7;bcd0<=5; end
			8576: begin bcd3<=8;bcd2<=5;bcd1<=7;bcd0<=6; end
			8577: begin bcd3<=8;bcd2<=5;bcd1<=7;bcd0<=7; end
			8578: begin bcd3<=8;bcd2<=5;bcd1<=7;bcd0<=8; end
			8579: begin bcd3<=8;bcd2<=5;bcd1<=7;bcd0<=9; end
			8580: begin bcd3<=8;bcd2<=5;bcd1<=8;bcd0<=0; end
			8581: begin bcd3<=8;bcd2<=5;bcd1<=8;bcd0<=1; end
			8582: begin bcd3<=8;bcd2<=5;bcd1<=8;bcd0<=2; end
			8583: begin bcd3<=8;bcd2<=5;bcd1<=8;bcd0<=3; end
			8584: begin bcd3<=8;bcd2<=5;bcd1<=8;bcd0<=4; end
			8585: begin bcd3<=8;bcd2<=5;bcd1<=8;bcd0<=5; end
			8586: begin bcd3<=8;bcd2<=5;bcd1<=8;bcd0<=6; end
			8587: begin bcd3<=8;bcd2<=5;bcd1<=8;bcd0<=7; end
			8588: begin bcd3<=8;bcd2<=5;bcd1<=8;bcd0<=8; end
			8589: begin bcd3<=8;bcd2<=5;bcd1<=8;bcd0<=9; end
			8590: begin bcd3<=8;bcd2<=5;bcd1<=9;bcd0<=0; end
			8591: begin bcd3<=8;bcd2<=5;bcd1<=9;bcd0<=1; end
			8592: begin bcd3<=8;bcd2<=5;bcd1<=9;bcd0<=2; end
			8593: begin bcd3<=8;bcd2<=5;bcd1<=9;bcd0<=3; end
			8594: begin bcd3<=8;bcd2<=5;bcd1<=9;bcd0<=4; end
			8595: begin bcd3<=8;bcd2<=5;bcd1<=9;bcd0<=5; end
			8596: begin bcd3<=8;bcd2<=5;bcd1<=9;bcd0<=6; end
			8597: begin bcd3<=8;bcd2<=5;bcd1<=9;bcd0<=7; end
			8598: begin bcd3<=8;bcd2<=5;bcd1<=9;bcd0<=8; end
			8599: begin bcd3<=8;bcd2<=5;bcd1<=9;bcd0<=9; end
			8600: begin bcd3<=8;bcd2<=6;bcd1<=0;bcd0<=0; end
			8601: begin bcd3<=8;bcd2<=6;bcd1<=0;bcd0<=1; end
			8602: begin bcd3<=8;bcd2<=6;bcd1<=0;bcd0<=2; end
			8603: begin bcd3<=8;bcd2<=6;bcd1<=0;bcd0<=3; end
			8604: begin bcd3<=8;bcd2<=6;bcd1<=0;bcd0<=4; end
			8605: begin bcd3<=8;bcd2<=6;bcd1<=0;bcd0<=5; end
			8606: begin bcd3<=8;bcd2<=6;bcd1<=0;bcd0<=6; end
			8607: begin bcd3<=8;bcd2<=6;bcd1<=0;bcd0<=7; end
			8608: begin bcd3<=8;bcd2<=6;bcd1<=0;bcd0<=8; end
			8609: begin bcd3<=8;bcd2<=6;bcd1<=0;bcd0<=9; end
			8610: begin bcd3<=8;bcd2<=6;bcd1<=1;bcd0<=0; end
			8611: begin bcd3<=8;bcd2<=6;bcd1<=1;bcd0<=1; end
			8612: begin bcd3<=8;bcd2<=6;bcd1<=1;bcd0<=2; end
			8613: begin bcd3<=8;bcd2<=6;bcd1<=1;bcd0<=3; end
			8614: begin bcd3<=8;bcd2<=6;bcd1<=1;bcd0<=4; end
			8615: begin bcd3<=8;bcd2<=6;bcd1<=1;bcd0<=5; end
			8616: begin bcd3<=8;bcd2<=6;bcd1<=1;bcd0<=6; end
			8617: begin bcd3<=8;bcd2<=6;bcd1<=1;bcd0<=7; end
			8618: begin bcd3<=8;bcd2<=6;bcd1<=1;bcd0<=8; end
			8619: begin bcd3<=8;bcd2<=6;bcd1<=1;bcd0<=9; end
			8620: begin bcd3<=8;bcd2<=6;bcd1<=2;bcd0<=0; end
			8621: begin bcd3<=8;bcd2<=6;bcd1<=2;bcd0<=1; end
			8622: begin bcd3<=8;bcd2<=6;bcd1<=2;bcd0<=2; end
			8623: begin bcd3<=8;bcd2<=6;bcd1<=2;bcd0<=3; end
			8624: begin bcd3<=8;bcd2<=6;bcd1<=2;bcd0<=4; end
			8625: begin bcd3<=8;bcd2<=6;bcd1<=2;bcd0<=5; end
			8626: begin bcd3<=8;bcd2<=6;bcd1<=2;bcd0<=6; end
			8627: begin bcd3<=8;bcd2<=6;bcd1<=2;bcd0<=7; end
			8628: begin bcd3<=8;bcd2<=6;bcd1<=2;bcd0<=8; end
			8629: begin bcd3<=8;bcd2<=6;bcd1<=2;bcd0<=9; end
			8630: begin bcd3<=8;bcd2<=6;bcd1<=3;bcd0<=0; end
			8631: begin bcd3<=8;bcd2<=6;bcd1<=3;bcd0<=1; end
			8632: begin bcd3<=8;bcd2<=6;bcd1<=3;bcd0<=2; end
			8633: begin bcd3<=8;bcd2<=6;bcd1<=3;bcd0<=3; end
			8634: begin bcd3<=8;bcd2<=6;bcd1<=3;bcd0<=4; end
			8635: begin bcd3<=8;bcd2<=6;bcd1<=3;bcd0<=5; end
			8636: begin bcd3<=8;bcd2<=6;bcd1<=3;bcd0<=6; end
			8637: begin bcd3<=8;bcd2<=6;bcd1<=3;bcd0<=7; end
			8638: begin bcd3<=8;bcd2<=6;bcd1<=3;bcd0<=8; end
			8639: begin bcd3<=8;bcd2<=6;bcd1<=3;bcd0<=9; end
			8640: begin bcd3<=8;bcd2<=6;bcd1<=4;bcd0<=0; end
			8641: begin bcd3<=8;bcd2<=6;bcd1<=4;bcd0<=1; end
			8642: begin bcd3<=8;bcd2<=6;bcd1<=4;bcd0<=2; end
			8643: begin bcd3<=8;bcd2<=6;bcd1<=4;bcd0<=3; end
			8644: begin bcd3<=8;bcd2<=6;bcd1<=4;bcd0<=4; end
			8645: begin bcd3<=8;bcd2<=6;bcd1<=4;bcd0<=5; end
			8646: begin bcd3<=8;bcd2<=6;bcd1<=4;bcd0<=6; end
			8647: begin bcd3<=8;bcd2<=6;bcd1<=4;bcd0<=7; end
			8648: begin bcd3<=8;bcd2<=6;bcd1<=4;bcd0<=8; end
			8649: begin bcd3<=8;bcd2<=6;bcd1<=4;bcd0<=9; end
			8650: begin bcd3<=8;bcd2<=6;bcd1<=5;bcd0<=0; end
			8651: begin bcd3<=8;bcd2<=6;bcd1<=5;bcd0<=1; end
			8652: begin bcd3<=8;bcd2<=6;bcd1<=5;bcd0<=2; end
			8653: begin bcd3<=8;bcd2<=6;bcd1<=5;bcd0<=3; end
			8654: begin bcd3<=8;bcd2<=6;bcd1<=5;bcd0<=4; end
			8655: begin bcd3<=8;bcd2<=6;bcd1<=5;bcd0<=5; end
			8656: begin bcd3<=8;bcd2<=6;bcd1<=5;bcd0<=6; end
			8657: begin bcd3<=8;bcd2<=6;bcd1<=5;bcd0<=7; end
			8658: begin bcd3<=8;bcd2<=6;bcd1<=5;bcd0<=8; end
			8659: begin bcd3<=8;bcd2<=6;bcd1<=5;bcd0<=9; end
			8660: begin bcd3<=8;bcd2<=6;bcd1<=6;bcd0<=0; end
			8661: begin bcd3<=8;bcd2<=6;bcd1<=6;bcd0<=1; end
			8662: begin bcd3<=8;bcd2<=6;bcd1<=6;bcd0<=2; end
			8663: begin bcd3<=8;bcd2<=6;bcd1<=6;bcd0<=3; end
			8664: begin bcd3<=8;bcd2<=6;bcd1<=6;bcd0<=4; end
			8665: begin bcd3<=8;bcd2<=6;bcd1<=6;bcd0<=5; end
			8666: begin bcd3<=8;bcd2<=6;bcd1<=6;bcd0<=6; end
			8667: begin bcd3<=8;bcd2<=6;bcd1<=6;bcd0<=7; end
			8668: begin bcd3<=8;bcd2<=6;bcd1<=6;bcd0<=8; end
			8669: begin bcd3<=8;bcd2<=6;bcd1<=6;bcd0<=9; end
			8670: begin bcd3<=8;bcd2<=6;bcd1<=7;bcd0<=0; end
			8671: begin bcd3<=8;bcd2<=6;bcd1<=7;bcd0<=1; end
			8672: begin bcd3<=8;bcd2<=6;bcd1<=7;bcd0<=2; end
			8673: begin bcd3<=8;bcd2<=6;bcd1<=7;bcd0<=3; end
			8674: begin bcd3<=8;bcd2<=6;bcd1<=7;bcd0<=4; end
			8675: begin bcd3<=8;bcd2<=6;bcd1<=7;bcd0<=5; end
			8676: begin bcd3<=8;bcd2<=6;bcd1<=7;bcd0<=6; end
			8677: begin bcd3<=8;bcd2<=6;bcd1<=7;bcd0<=7; end
			8678: begin bcd3<=8;bcd2<=6;bcd1<=7;bcd0<=8; end
			8679: begin bcd3<=8;bcd2<=6;bcd1<=7;bcd0<=9; end
			8680: begin bcd3<=8;bcd2<=6;bcd1<=8;bcd0<=0; end
			8681: begin bcd3<=8;bcd2<=6;bcd1<=8;bcd0<=1; end
			8682: begin bcd3<=8;bcd2<=6;bcd1<=8;bcd0<=2; end
			8683: begin bcd3<=8;bcd2<=6;bcd1<=8;bcd0<=3; end
			8684: begin bcd3<=8;bcd2<=6;bcd1<=8;bcd0<=4; end
			8685: begin bcd3<=8;bcd2<=6;bcd1<=8;bcd0<=5; end
			8686: begin bcd3<=8;bcd2<=6;bcd1<=8;bcd0<=6; end
			8687: begin bcd3<=8;bcd2<=6;bcd1<=8;bcd0<=7; end
			8688: begin bcd3<=8;bcd2<=6;bcd1<=8;bcd0<=8; end
			8689: begin bcd3<=8;bcd2<=6;bcd1<=8;bcd0<=9; end
			8690: begin bcd3<=8;bcd2<=6;bcd1<=9;bcd0<=0; end
			8691: begin bcd3<=8;bcd2<=6;bcd1<=9;bcd0<=1; end
			8692: begin bcd3<=8;bcd2<=6;bcd1<=9;bcd0<=2; end
			8693: begin bcd3<=8;bcd2<=6;bcd1<=9;bcd0<=3; end
			8694: begin bcd3<=8;bcd2<=6;bcd1<=9;bcd0<=4; end
			8695: begin bcd3<=8;bcd2<=6;bcd1<=9;bcd0<=5; end
			8696: begin bcd3<=8;bcd2<=6;bcd1<=9;bcd0<=6; end
			8697: begin bcd3<=8;bcd2<=6;bcd1<=9;bcd0<=7; end
			8698: begin bcd3<=8;bcd2<=6;bcd1<=9;bcd0<=8; end
			8699: begin bcd3<=8;bcd2<=6;bcd1<=9;bcd0<=9; end
			8700: begin bcd3<=8;bcd2<=7;bcd1<=0;bcd0<=0; end
			8701: begin bcd3<=8;bcd2<=7;bcd1<=0;bcd0<=1; end
			8702: begin bcd3<=8;bcd2<=7;bcd1<=0;bcd0<=2; end
			8703: begin bcd3<=8;bcd2<=7;bcd1<=0;bcd0<=3; end
			8704: begin bcd3<=8;bcd2<=7;bcd1<=0;bcd0<=4; end
			8705: begin bcd3<=8;bcd2<=7;bcd1<=0;bcd0<=5; end
			8706: begin bcd3<=8;bcd2<=7;bcd1<=0;bcd0<=6; end
			8707: begin bcd3<=8;bcd2<=7;bcd1<=0;bcd0<=7; end
			8708: begin bcd3<=8;bcd2<=7;bcd1<=0;bcd0<=8; end
			8709: begin bcd3<=8;bcd2<=7;bcd1<=0;bcd0<=9; end
			8710: begin bcd3<=8;bcd2<=7;bcd1<=1;bcd0<=0; end
			8711: begin bcd3<=8;bcd2<=7;bcd1<=1;bcd0<=1; end
			8712: begin bcd3<=8;bcd2<=7;bcd1<=1;bcd0<=2; end
			8713: begin bcd3<=8;bcd2<=7;bcd1<=1;bcd0<=3; end
			8714: begin bcd3<=8;bcd2<=7;bcd1<=1;bcd0<=4; end
			8715: begin bcd3<=8;bcd2<=7;bcd1<=1;bcd0<=5; end
			8716: begin bcd3<=8;bcd2<=7;bcd1<=1;bcd0<=6; end
			8717: begin bcd3<=8;bcd2<=7;bcd1<=1;bcd0<=7; end
			8718: begin bcd3<=8;bcd2<=7;bcd1<=1;bcd0<=8; end
			8719: begin bcd3<=8;bcd2<=7;bcd1<=1;bcd0<=9; end
			8720: begin bcd3<=8;bcd2<=7;bcd1<=2;bcd0<=0; end
			8721: begin bcd3<=8;bcd2<=7;bcd1<=2;bcd0<=1; end
			8722: begin bcd3<=8;bcd2<=7;bcd1<=2;bcd0<=2; end
			8723: begin bcd3<=8;bcd2<=7;bcd1<=2;bcd0<=3; end
			8724: begin bcd3<=8;bcd2<=7;bcd1<=2;bcd0<=4; end
			8725: begin bcd3<=8;bcd2<=7;bcd1<=2;bcd0<=5; end
			8726: begin bcd3<=8;bcd2<=7;bcd1<=2;bcd0<=6; end
			8727: begin bcd3<=8;bcd2<=7;bcd1<=2;bcd0<=7; end
			8728: begin bcd3<=8;bcd2<=7;bcd1<=2;bcd0<=8; end
			8729: begin bcd3<=8;bcd2<=7;bcd1<=2;bcd0<=9; end
			8730: begin bcd3<=8;bcd2<=7;bcd1<=3;bcd0<=0; end
			8731: begin bcd3<=8;bcd2<=7;bcd1<=3;bcd0<=1; end
			8732: begin bcd3<=8;bcd2<=7;bcd1<=3;bcd0<=2; end
			8733: begin bcd3<=8;bcd2<=7;bcd1<=3;bcd0<=3; end
			8734: begin bcd3<=8;bcd2<=7;bcd1<=3;bcd0<=4; end
			8735: begin bcd3<=8;bcd2<=7;bcd1<=3;bcd0<=5; end
			8736: begin bcd3<=8;bcd2<=7;bcd1<=3;bcd0<=6; end
			8737: begin bcd3<=8;bcd2<=7;bcd1<=3;bcd0<=7; end
			8738: begin bcd3<=8;bcd2<=7;bcd1<=3;bcd0<=8; end
			8739: begin bcd3<=8;bcd2<=7;bcd1<=3;bcd0<=9; end
			8740: begin bcd3<=8;bcd2<=7;bcd1<=4;bcd0<=0; end
			8741: begin bcd3<=8;bcd2<=7;bcd1<=4;bcd0<=1; end
			8742: begin bcd3<=8;bcd2<=7;bcd1<=4;bcd0<=2; end
			8743: begin bcd3<=8;bcd2<=7;bcd1<=4;bcd0<=3; end
			8744: begin bcd3<=8;bcd2<=7;bcd1<=4;bcd0<=4; end
			8745: begin bcd3<=8;bcd2<=7;bcd1<=4;bcd0<=5; end
			8746: begin bcd3<=8;bcd2<=7;bcd1<=4;bcd0<=6; end
			8747: begin bcd3<=8;bcd2<=7;bcd1<=4;bcd0<=7; end
			8748: begin bcd3<=8;bcd2<=7;bcd1<=4;bcd0<=8; end
			8749: begin bcd3<=8;bcd2<=7;bcd1<=4;bcd0<=9; end
			8750: begin bcd3<=8;bcd2<=7;bcd1<=5;bcd0<=0; end
			8751: begin bcd3<=8;bcd2<=7;bcd1<=5;bcd0<=1; end
			8752: begin bcd3<=8;bcd2<=7;bcd1<=5;bcd0<=2; end
			8753: begin bcd3<=8;bcd2<=7;bcd1<=5;bcd0<=3; end
			8754: begin bcd3<=8;bcd2<=7;bcd1<=5;bcd0<=4; end
			8755: begin bcd3<=8;bcd2<=7;bcd1<=5;bcd0<=5; end
			8756: begin bcd3<=8;bcd2<=7;bcd1<=5;bcd0<=6; end
			8757: begin bcd3<=8;bcd2<=7;bcd1<=5;bcd0<=7; end
			8758: begin bcd3<=8;bcd2<=7;bcd1<=5;bcd0<=8; end
			8759: begin bcd3<=8;bcd2<=7;bcd1<=5;bcd0<=9; end
			8760: begin bcd3<=8;bcd2<=7;bcd1<=6;bcd0<=0; end
			8761: begin bcd3<=8;bcd2<=7;bcd1<=6;bcd0<=1; end
			8762: begin bcd3<=8;bcd2<=7;bcd1<=6;bcd0<=2; end
			8763: begin bcd3<=8;bcd2<=7;bcd1<=6;bcd0<=3; end
			8764: begin bcd3<=8;bcd2<=7;bcd1<=6;bcd0<=4; end
			8765: begin bcd3<=8;bcd2<=7;bcd1<=6;bcd0<=5; end
			8766: begin bcd3<=8;bcd2<=7;bcd1<=6;bcd0<=6; end
			8767: begin bcd3<=8;bcd2<=7;bcd1<=6;bcd0<=7; end
			8768: begin bcd3<=8;bcd2<=7;bcd1<=6;bcd0<=8; end
			8769: begin bcd3<=8;bcd2<=7;bcd1<=6;bcd0<=9; end
			8770: begin bcd3<=8;bcd2<=7;bcd1<=7;bcd0<=0; end
			8771: begin bcd3<=8;bcd2<=7;bcd1<=7;bcd0<=1; end
			8772: begin bcd3<=8;bcd2<=7;bcd1<=7;bcd0<=2; end
			8773: begin bcd3<=8;bcd2<=7;bcd1<=7;bcd0<=3; end
			8774: begin bcd3<=8;bcd2<=7;bcd1<=7;bcd0<=4; end
			8775: begin bcd3<=8;bcd2<=7;bcd1<=7;bcd0<=5; end
			8776: begin bcd3<=8;bcd2<=7;bcd1<=7;bcd0<=6; end
			8777: begin bcd3<=8;bcd2<=7;bcd1<=7;bcd0<=7; end
			8778: begin bcd3<=8;bcd2<=7;bcd1<=7;bcd0<=8; end
			8779: begin bcd3<=8;bcd2<=7;bcd1<=7;bcd0<=9; end
			8780: begin bcd3<=8;bcd2<=7;bcd1<=8;bcd0<=0; end
			8781: begin bcd3<=8;bcd2<=7;bcd1<=8;bcd0<=1; end
			8782: begin bcd3<=8;bcd2<=7;bcd1<=8;bcd0<=2; end
			8783: begin bcd3<=8;bcd2<=7;bcd1<=8;bcd0<=3; end
			8784: begin bcd3<=8;bcd2<=7;bcd1<=8;bcd0<=4; end
			8785: begin bcd3<=8;bcd2<=7;bcd1<=8;bcd0<=5; end
			8786: begin bcd3<=8;bcd2<=7;bcd1<=8;bcd0<=6; end
			8787: begin bcd3<=8;bcd2<=7;bcd1<=8;bcd0<=7; end
			8788: begin bcd3<=8;bcd2<=7;bcd1<=8;bcd0<=8; end
			8789: begin bcd3<=8;bcd2<=7;bcd1<=8;bcd0<=9; end
			8790: begin bcd3<=8;bcd2<=7;bcd1<=9;bcd0<=0; end
			8791: begin bcd3<=8;bcd2<=7;bcd1<=9;bcd0<=1; end
			8792: begin bcd3<=8;bcd2<=7;bcd1<=9;bcd0<=2; end
			8793: begin bcd3<=8;bcd2<=7;bcd1<=9;bcd0<=3; end
			8794: begin bcd3<=8;bcd2<=7;bcd1<=9;bcd0<=4; end
			8795: begin bcd3<=8;bcd2<=7;bcd1<=9;bcd0<=5; end
			8796: begin bcd3<=8;bcd2<=7;bcd1<=9;bcd0<=6; end
			8797: begin bcd3<=8;bcd2<=7;bcd1<=9;bcd0<=7; end
			8798: begin bcd3<=8;bcd2<=7;bcd1<=9;bcd0<=8; end
			8799: begin bcd3<=8;bcd2<=7;bcd1<=9;bcd0<=9; end
			8800: begin bcd3<=8;bcd2<=8;bcd1<=0;bcd0<=0; end
			8801: begin bcd3<=8;bcd2<=8;bcd1<=0;bcd0<=1; end
			8802: begin bcd3<=8;bcd2<=8;bcd1<=0;bcd0<=2; end
			8803: begin bcd3<=8;bcd2<=8;bcd1<=0;bcd0<=3; end
			8804: begin bcd3<=8;bcd2<=8;bcd1<=0;bcd0<=4; end
			8805: begin bcd3<=8;bcd2<=8;bcd1<=0;bcd0<=5; end
			8806: begin bcd3<=8;bcd2<=8;bcd1<=0;bcd0<=6; end
			8807: begin bcd3<=8;bcd2<=8;bcd1<=0;bcd0<=7; end
			8808: begin bcd3<=8;bcd2<=8;bcd1<=0;bcd0<=8; end
			8809: begin bcd3<=8;bcd2<=8;bcd1<=0;bcd0<=9; end
			8810: begin bcd3<=8;bcd2<=8;bcd1<=1;bcd0<=0; end
			8811: begin bcd3<=8;bcd2<=8;bcd1<=1;bcd0<=1; end
			8812: begin bcd3<=8;bcd2<=8;bcd1<=1;bcd0<=2; end
			8813: begin bcd3<=8;bcd2<=8;bcd1<=1;bcd0<=3; end
			8814: begin bcd3<=8;bcd2<=8;bcd1<=1;bcd0<=4; end
			8815: begin bcd3<=8;bcd2<=8;bcd1<=1;bcd0<=5; end
			8816: begin bcd3<=8;bcd2<=8;bcd1<=1;bcd0<=6; end
			8817: begin bcd3<=8;bcd2<=8;bcd1<=1;bcd0<=7; end
			8818: begin bcd3<=8;bcd2<=8;bcd1<=1;bcd0<=8; end
			8819: begin bcd3<=8;bcd2<=8;bcd1<=1;bcd0<=9; end
			8820: begin bcd3<=8;bcd2<=8;bcd1<=2;bcd0<=0; end
			8821: begin bcd3<=8;bcd2<=8;bcd1<=2;bcd0<=1; end
			8822: begin bcd3<=8;bcd2<=8;bcd1<=2;bcd0<=2; end
			8823: begin bcd3<=8;bcd2<=8;bcd1<=2;bcd0<=3; end
			8824: begin bcd3<=8;bcd2<=8;bcd1<=2;bcd0<=4; end
			8825: begin bcd3<=8;bcd2<=8;bcd1<=2;bcd0<=5; end
			8826: begin bcd3<=8;bcd2<=8;bcd1<=2;bcd0<=6; end
			8827: begin bcd3<=8;bcd2<=8;bcd1<=2;bcd0<=7; end
			8828: begin bcd3<=8;bcd2<=8;bcd1<=2;bcd0<=8; end
			8829: begin bcd3<=8;bcd2<=8;bcd1<=2;bcd0<=9; end
			8830: begin bcd3<=8;bcd2<=8;bcd1<=3;bcd0<=0; end
			8831: begin bcd3<=8;bcd2<=8;bcd1<=3;bcd0<=1; end
			8832: begin bcd3<=8;bcd2<=8;bcd1<=3;bcd0<=2; end
			8833: begin bcd3<=8;bcd2<=8;bcd1<=3;bcd0<=3; end
			8834: begin bcd3<=8;bcd2<=8;bcd1<=3;bcd0<=4; end
			8835: begin bcd3<=8;bcd2<=8;bcd1<=3;bcd0<=5; end
			8836: begin bcd3<=8;bcd2<=8;bcd1<=3;bcd0<=6; end
			8837: begin bcd3<=8;bcd2<=8;bcd1<=3;bcd0<=7; end
			8838: begin bcd3<=8;bcd2<=8;bcd1<=3;bcd0<=8; end
			8839: begin bcd3<=8;bcd2<=8;bcd1<=3;bcd0<=9; end
			8840: begin bcd3<=8;bcd2<=8;bcd1<=4;bcd0<=0; end
			8841: begin bcd3<=8;bcd2<=8;bcd1<=4;bcd0<=1; end
			8842: begin bcd3<=8;bcd2<=8;bcd1<=4;bcd0<=2; end
			8843: begin bcd3<=8;bcd2<=8;bcd1<=4;bcd0<=3; end
			8844: begin bcd3<=8;bcd2<=8;bcd1<=4;bcd0<=4; end
			8845: begin bcd3<=8;bcd2<=8;bcd1<=4;bcd0<=5; end
			8846: begin bcd3<=8;bcd2<=8;bcd1<=4;bcd0<=6; end
			8847: begin bcd3<=8;bcd2<=8;bcd1<=4;bcd0<=7; end
			8848: begin bcd3<=8;bcd2<=8;bcd1<=4;bcd0<=8; end
			8849: begin bcd3<=8;bcd2<=8;bcd1<=4;bcd0<=9; end
			8850: begin bcd3<=8;bcd2<=8;bcd1<=5;bcd0<=0; end
			8851: begin bcd3<=8;bcd2<=8;bcd1<=5;bcd0<=1; end
			8852: begin bcd3<=8;bcd2<=8;bcd1<=5;bcd0<=2; end
			8853: begin bcd3<=8;bcd2<=8;bcd1<=5;bcd0<=3; end
			8854: begin bcd3<=8;bcd2<=8;bcd1<=5;bcd0<=4; end
			8855: begin bcd3<=8;bcd2<=8;bcd1<=5;bcd0<=5; end
			8856: begin bcd3<=8;bcd2<=8;bcd1<=5;bcd0<=6; end
			8857: begin bcd3<=8;bcd2<=8;bcd1<=5;bcd0<=7; end
			8858: begin bcd3<=8;bcd2<=8;bcd1<=5;bcd0<=8; end
			8859: begin bcd3<=8;bcd2<=8;bcd1<=5;bcd0<=9; end
			8860: begin bcd3<=8;bcd2<=8;bcd1<=6;bcd0<=0; end
			8861: begin bcd3<=8;bcd2<=8;bcd1<=6;bcd0<=1; end
			8862: begin bcd3<=8;bcd2<=8;bcd1<=6;bcd0<=2; end
			8863: begin bcd3<=8;bcd2<=8;bcd1<=6;bcd0<=3; end
			8864: begin bcd3<=8;bcd2<=8;bcd1<=6;bcd0<=4; end
			8865: begin bcd3<=8;bcd2<=8;bcd1<=6;bcd0<=5; end
			8866: begin bcd3<=8;bcd2<=8;bcd1<=6;bcd0<=6; end
			8867: begin bcd3<=8;bcd2<=8;bcd1<=6;bcd0<=7; end
			8868: begin bcd3<=8;bcd2<=8;bcd1<=6;bcd0<=8; end
			8869: begin bcd3<=8;bcd2<=8;bcd1<=6;bcd0<=9; end
			8870: begin bcd3<=8;bcd2<=8;bcd1<=7;bcd0<=0; end
			8871: begin bcd3<=8;bcd2<=8;bcd1<=7;bcd0<=1; end
			8872: begin bcd3<=8;bcd2<=8;bcd1<=7;bcd0<=2; end
			8873: begin bcd3<=8;bcd2<=8;bcd1<=7;bcd0<=3; end
			8874: begin bcd3<=8;bcd2<=8;bcd1<=7;bcd0<=4; end
			8875: begin bcd3<=8;bcd2<=8;bcd1<=7;bcd0<=5; end
			8876: begin bcd3<=8;bcd2<=8;bcd1<=7;bcd0<=6; end
			8877: begin bcd3<=8;bcd2<=8;bcd1<=7;bcd0<=7; end
			8878: begin bcd3<=8;bcd2<=8;bcd1<=7;bcd0<=8; end
			8879: begin bcd3<=8;bcd2<=8;bcd1<=7;bcd0<=9; end
			8880: begin bcd3<=8;bcd2<=8;bcd1<=8;bcd0<=0; end
			8881: begin bcd3<=8;bcd2<=8;bcd1<=8;bcd0<=1; end
			8882: begin bcd3<=8;bcd2<=8;bcd1<=8;bcd0<=2; end
			8883: begin bcd3<=8;bcd2<=8;bcd1<=8;bcd0<=3; end
			8884: begin bcd3<=8;bcd2<=8;bcd1<=8;bcd0<=4; end
			8885: begin bcd3<=8;bcd2<=8;bcd1<=8;bcd0<=5; end
			8886: begin bcd3<=8;bcd2<=8;bcd1<=8;bcd0<=6; end
			8887: begin bcd3<=8;bcd2<=8;bcd1<=8;bcd0<=7; end
			8888: begin bcd3<=8;bcd2<=8;bcd1<=8;bcd0<=8; end
			8889: begin bcd3<=8;bcd2<=8;bcd1<=8;bcd0<=9; end
			8890: begin bcd3<=8;bcd2<=8;bcd1<=9;bcd0<=0; end
			8891: begin bcd3<=8;bcd2<=8;bcd1<=9;bcd0<=1; end
			8892: begin bcd3<=8;bcd2<=8;bcd1<=9;bcd0<=2; end
			8893: begin bcd3<=8;bcd2<=8;bcd1<=9;bcd0<=3; end
			8894: begin bcd3<=8;bcd2<=8;bcd1<=9;bcd0<=4; end
			8895: begin bcd3<=8;bcd2<=8;bcd1<=9;bcd0<=5; end
			8896: begin bcd3<=8;bcd2<=8;bcd1<=9;bcd0<=6; end
			8897: begin bcd3<=8;bcd2<=8;bcd1<=9;bcd0<=7; end
			8898: begin bcd3<=8;bcd2<=8;bcd1<=9;bcd0<=8; end
			8899: begin bcd3<=8;bcd2<=8;bcd1<=9;bcd0<=9; end
			8900: begin bcd3<=8;bcd2<=9;bcd1<=0;bcd0<=0; end
			8901: begin bcd3<=8;bcd2<=9;bcd1<=0;bcd0<=1; end
			8902: begin bcd3<=8;bcd2<=9;bcd1<=0;bcd0<=2; end
			8903: begin bcd3<=8;bcd2<=9;bcd1<=0;bcd0<=3; end
			8904: begin bcd3<=8;bcd2<=9;bcd1<=0;bcd0<=4; end
			8905: begin bcd3<=8;bcd2<=9;bcd1<=0;bcd0<=5; end
			8906: begin bcd3<=8;bcd2<=9;bcd1<=0;bcd0<=6; end
			8907: begin bcd3<=8;bcd2<=9;bcd1<=0;bcd0<=7; end
			8908: begin bcd3<=8;bcd2<=9;bcd1<=0;bcd0<=8; end
			8909: begin bcd3<=8;bcd2<=9;bcd1<=0;bcd0<=9; end
			8910: begin bcd3<=8;bcd2<=9;bcd1<=1;bcd0<=0; end
			8911: begin bcd3<=8;bcd2<=9;bcd1<=1;bcd0<=1; end
			8912: begin bcd3<=8;bcd2<=9;bcd1<=1;bcd0<=2; end
			8913: begin bcd3<=8;bcd2<=9;bcd1<=1;bcd0<=3; end
			8914: begin bcd3<=8;bcd2<=9;bcd1<=1;bcd0<=4; end
			8915: begin bcd3<=8;bcd2<=9;bcd1<=1;bcd0<=5; end
			8916: begin bcd3<=8;bcd2<=9;bcd1<=1;bcd0<=6; end
			8917: begin bcd3<=8;bcd2<=9;bcd1<=1;bcd0<=7; end
			8918: begin bcd3<=8;bcd2<=9;bcd1<=1;bcd0<=8; end
			8919: begin bcd3<=8;bcd2<=9;bcd1<=1;bcd0<=9; end
			8920: begin bcd3<=8;bcd2<=9;bcd1<=2;bcd0<=0; end
			8921: begin bcd3<=8;bcd2<=9;bcd1<=2;bcd0<=1; end
			8922: begin bcd3<=8;bcd2<=9;bcd1<=2;bcd0<=2; end
			8923: begin bcd3<=8;bcd2<=9;bcd1<=2;bcd0<=3; end
			8924: begin bcd3<=8;bcd2<=9;bcd1<=2;bcd0<=4; end
			8925: begin bcd3<=8;bcd2<=9;bcd1<=2;bcd0<=5; end
			8926: begin bcd3<=8;bcd2<=9;bcd1<=2;bcd0<=6; end
			8927: begin bcd3<=8;bcd2<=9;bcd1<=2;bcd0<=7; end
			8928: begin bcd3<=8;bcd2<=9;bcd1<=2;bcd0<=8; end
			8929: begin bcd3<=8;bcd2<=9;bcd1<=2;bcd0<=9; end
			8930: begin bcd3<=8;bcd2<=9;bcd1<=3;bcd0<=0; end
			8931: begin bcd3<=8;bcd2<=9;bcd1<=3;bcd0<=1; end
			8932: begin bcd3<=8;bcd2<=9;bcd1<=3;bcd0<=2; end
			8933: begin bcd3<=8;bcd2<=9;bcd1<=3;bcd0<=3; end
			8934: begin bcd3<=8;bcd2<=9;bcd1<=3;bcd0<=4; end
			8935: begin bcd3<=8;bcd2<=9;bcd1<=3;bcd0<=5; end
			8936: begin bcd3<=8;bcd2<=9;bcd1<=3;bcd0<=6; end
			8937: begin bcd3<=8;bcd2<=9;bcd1<=3;bcd0<=7; end
			8938: begin bcd3<=8;bcd2<=9;bcd1<=3;bcd0<=8; end
			8939: begin bcd3<=8;bcd2<=9;bcd1<=3;bcd0<=9; end
			8940: begin bcd3<=8;bcd2<=9;bcd1<=4;bcd0<=0; end
			8941: begin bcd3<=8;bcd2<=9;bcd1<=4;bcd0<=1; end
			8942: begin bcd3<=8;bcd2<=9;bcd1<=4;bcd0<=2; end
			8943: begin bcd3<=8;bcd2<=9;bcd1<=4;bcd0<=3; end
			8944: begin bcd3<=8;bcd2<=9;bcd1<=4;bcd0<=4; end
			8945: begin bcd3<=8;bcd2<=9;bcd1<=4;bcd0<=5; end
			8946: begin bcd3<=8;bcd2<=9;bcd1<=4;bcd0<=6; end
			8947: begin bcd3<=8;bcd2<=9;bcd1<=4;bcd0<=7; end
			8948: begin bcd3<=8;bcd2<=9;bcd1<=4;bcd0<=8; end
			8949: begin bcd3<=8;bcd2<=9;bcd1<=4;bcd0<=9; end
			8950: begin bcd3<=8;bcd2<=9;bcd1<=5;bcd0<=0; end
			8951: begin bcd3<=8;bcd2<=9;bcd1<=5;bcd0<=1; end
			8952: begin bcd3<=8;bcd2<=9;bcd1<=5;bcd0<=2; end
			8953: begin bcd3<=8;bcd2<=9;bcd1<=5;bcd0<=3; end
			8954: begin bcd3<=8;bcd2<=9;bcd1<=5;bcd0<=4; end
			8955: begin bcd3<=8;bcd2<=9;bcd1<=5;bcd0<=5; end
			8956: begin bcd3<=8;bcd2<=9;bcd1<=5;bcd0<=6; end
			8957: begin bcd3<=8;bcd2<=9;bcd1<=5;bcd0<=7; end
			8958: begin bcd3<=8;bcd2<=9;bcd1<=5;bcd0<=8; end
			8959: begin bcd3<=8;bcd2<=9;bcd1<=5;bcd0<=9; end
			8960: begin bcd3<=8;bcd2<=9;bcd1<=6;bcd0<=0; end
			8961: begin bcd3<=8;bcd2<=9;bcd1<=6;bcd0<=1; end
			8962: begin bcd3<=8;bcd2<=9;bcd1<=6;bcd0<=2; end
			8963: begin bcd3<=8;bcd2<=9;bcd1<=6;bcd0<=3; end
			8964: begin bcd3<=8;bcd2<=9;bcd1<=6;bcd0<=4; end
			8965: begin bcd3<=8;bcd2<=9;bcd1<=6;bcd0<=5; end
			8966: begin bcd3<=8;bcd2<=9;bcd1<=6;bcd0<=6; end
			8967: begin bcd3<=8;bcd2<=9;bcd1<=6;bcd0<=7; end
			8968: begin bcd3<=8;bcd2<=9;bcd1<=6;bcd0<=8; end
			8969: begin bcd3<=8;bcd2<=9;bcd1<=6;bcd0<=9; end
			8970: begin bcd3<=8;bcd2<=9;bcd1<=7;bcd0<=0; end
			8971: begin bcd3<=8;bcd2<=9;bcd1<=7;bcd0<=1; end
			8972: begin bcd3<=8;bcd2<=9;bcd1<=7;bcd0<=2; end
			8973: begin bcd3<=8;bcd2<=9;bcd1<=7;bcd0<=3; end
			8974: begin bcd3<=8;bcd2<=9;bcd1<=7;bcd0<=4; end
			8975: begin bcd3<=8;bcd2<=9;bcd1<=7;bcd0<=5; end
			8976: begin bcd3<=8;bcd2<=9;bcd1<=7;bcd0<=6; end
			8977: begin bcd3<=8;bcd2<=9;bcd1<=7;bcd0<=7; end
			8978: begin bcd3<=8;bcd2<=9;bcd1<=7;bcd0<=8; end
			8979: begin bcd3<=8;bcd2<=9;bcd1<=7;bcd0<=9; end
			8980: begin bcd3<=8;bcd2<=9;bcd1<=8;bcd0<=0; end
			8981: begin bcd3<=8;bcd2<=9;bcd1<=8;bcd0<=1; end
			8982: begin bcd3<=8;bcd2<=9;bcd1<=8;bcd0<=2; end
			8983: begin bcd3<=8;bcd2<=9;bcd1<=8;bcd0<=3; end
			8984: begin bcd3<=8;bcd2<=9;bcd1<=8;bcd0<=4; end
			8985: begin bcd3<=8;bcd2<=9;bcd1<=8;bcd0<=5; end
			8986: begin bcd3<=8;bcd2<=9;bcd1<=8;bcd0<=6; end
			8987: begin bcd3<=8;bcd2<=9;bcd1<=8;bcd0<=7; end
			8988: begin bcd3<=8;bcd2<=9;bcd1<=8;bcd0<=8; end
			8989: begin bcd3<=8;bcd2<=9;bcd1<=8;bcd0<=9; end
			8990: begin bcd3<=8;bcd2<=9;bcd1<=9;bcd0<=0; end
			8991: begin bcd3<=8;bcd2<=9;bcd1<=9;bcd0<=1; end
			8992: begin bcd3<=8;bcd2<=9;bcd1<=9;bcd0<=2; end
			8993: begin bcd3<=8;bcd2<=9;bcd1<=9;bcd0<=3; end
			8994: begin bcd3<=8;bcd2<=9;bcd1<=9;bcd0<=4; end
			8995: begin bcd3<=8;bcd2<=9;bcd1<=9;bcd0<=5; end
			8996: begin bcd3<=8;bcd2<=9;bcd1<=9;bcd0<=6; end
			8997: begin bcd3<=8;bcd2<=9;bcd1<=9;bcd0<=7; end
			8998: begin bcd3<=8;bcd2<=9;bcd1<=9;bcd0<=8; end
			8999: begin bcd3<=8;bcd2<=9;bcd1<=9;bcd0<=9; end
			9000: begin bcd3<=9;bcd2<=0;bcd1<=0;bcd0<=0; end
			9001: begin bcd3<=9;bcd2<=0;bcd1<=0;bcd0<=1; end
			9002: begin bcd3<=9;bcd2<=0;bcd1<=0;bcd0<=2; end
			9003: begin bcd3<=9;bcd2<=0;bcd1<=0;bcd0<=3; end
			9004: begin bcd3<=9;bcd2<=0;bcd1<=0;bcd0<=4; end
			9005: begin bcd3<=9;bcd2<=0;bcd1<=0;bcd0<=5; end
			9006: begin bcd3<=9;bcd2<=0;bcd1<=0;bcd0<=6; end
			9007: begin bcd3<=9;bcd2<=0;bcd1<=0;bcd0<=7; end
			9008: begin bcd3<=9;bcd2<=0;bcd1<=0;bcd0<=8; end
			9009: begin bcd3<=9;bcd2<=0;bcd1<=0;bcd0<=9; end
			9010: begin bcd3<=9;bcd2<=0;bcd1<=1;bcd0<=0; end
			9011: begin bcd3<=9;bcd2<=0;bcd1<=1;bcd0<=1; end
			9012: begin bcd3<=9;bcd2<=0;bcd1<=1;bcd0<=2; end
			9013: begin bcd3<=9;bcd2<=0;bcd1<=1;bcd0<=3; end
			9014: begin bcd3<=9;bcd2<=0;bcd1<=1;bcd0<=4; end
			9015: begin bcd3<=9;bcd2<=0;bcd1<=1;bcd0<=5; end
			9016: begin bcd3<=9;bcd2<=0;bcd1<=1;bcd0<=6; end
			9017: begin bcd3<=9;bcd2<=0;bcd1<=1;bcd0<=7; end
			9018: begin bcd3<=9;bcd2<=0;bcd1<=1;bcd0<=8; end
			9019: begin bcd3<=9;bcd2<=0;bcd1<=1;bcd0<=9; end
			9020: begin bcd3<=9;bcd2<=0;bcd1<=2;bcd0<=0; end
			9021: begin bcd3<=9;bcd2<=0;bcd1<=2;bcd0<=1; end
			9022: begin bcd3<=9;bcd2<=0;bcd1<=2;bcd0<=2; end
			9023: begin bcd3<=9;bcd2<=0;bcd1<=2;bcd0<=3; end
			9024: begin bcd3<=9;bcd2<=0;bcd1<=2;bcd0<=4; end
			9025: begin bcd3<=9;bcd2<=0;bcd1<=2;bcd0<=5; end
			9026: begin bcd3<=9;bcd2<=0;bcd1<=2;bcd0<=6; end
			9027: begin bcd3<=9;bcd2<=0;bcd1<=2;bcd0<=7; end
			9028: begin bcd3<=9;bcd2<=0;bcd1<=2;bcd0<=8; end
			9029: begin bcd3<=9;bcd2<=0;bcd1<=2;bcd0<=9; end
			9030: begin bcd3<=9;bcd2<=0;bcd1<=3;bcd0<=0; end
			9031: begin bcd3<=9;bcd2<=0;bcd1<=3;bcd0<=1; end
			9032: begin bcd3<=9;bcd2<=0;bcd1<=3;bcd0<=2; end
			9033: begin bcd3<=9;bcd2<=0;bcd1<=3;bcd0<=3; end
			9034: begin bcd3<=9;bcd2<=0;bcd1<=3;bcd0<=4; end
			9035: begin bcd3<=9;bcd2<=0;bcd1<=3;bcd0<=5; end
			9036: begin bcd3<=9;bcd2<=0;bcd1<=3;bcd0<=6; end
			9037: begin bcd3<=9;bcd2<=0;bcd1<=3;bcd0<=7; end
			9038: begin bcd3<=9;bcd2<=0;bcd1<=3;bcd0<=8; end
			9039: begin bcd3<=9;bcd2<=0;bcd1<=3;bcd0<=9; end
			9040: begin bcd3<=9;bcd2<=0;bcd1<=4;bcd0<=0; end
			9041: begin bcd3<=9;bcd2<=0;bcd1<=4;bcd0<=1; end
			9042: begin bcd3<=9;bcd2<=0;bcd1<=4;bcd0<=2; end
			9043: begin bcd3<=9;bcd2<=0;bcd1<=4;bcd0<=3; end
			9044: begin bcd3<=9;bcd2<=0;bcd1<=4;bcd0<=4; end
			9045: begin bcd3<=9;bcd2<=0;bcd1<=4;bcd0<=5; end
			9046: begin bcd3<=9;bcd2<=0;bcd1<=4;bcd0<=6; end
			9047: begin bcd3<=9;bcd2<=0;bcd1<=4;bcd0<=7; end
			9048: begin bcd3<=9;bcd2<=0;bcd1<=4;bcd0<=8; end
			9049: begin bcd3<=9;bcd2<=0;bcd1<=4;bcd0<=9; end
			9050: begin bcd3<=9;bcd2<=0;bcd1<=5;bcd0<=0; end
			9051: begin bcd3<=9;bcd2<=0;bcd1<=5;bcd0<=1; end
			9052: begin bcd3<=9;bcd2<=0;bcd1<=5;bcd0<=2; end
			9053: begin bcd3<=9;bcd2<=0;bcd1<=5;bcd0<=3; end
			9054: begin bcd3<=9;bcd2<=0;bcd1<=5;bcd0<=4; end
			9055: begin bcd3<=9;bcd2<=0;bcd1<=5;bcd0<=5; end
			9056: begin bcd3<=9;bcd2<=0;bcd1<=5;bcd0<=6; end
			9057: begin bcd3<=9;bcd2<=0;bcd1<=5;bcd0<=7; end
			9058: begin bcd3<=9;bcd2<=0;bcd1<=5;bcd0<=8; end
			9059: begin bcd3<=9;bcd2<=0;bcd1<=5;bcd0<=9; end
			9060: begin bcd3<=9;bcd2<=0;bcd1<=6;bcd0<=0; end
			9061: begin bcd3<=9;bcd2<=0;bcd1<=6;bcd0<=1; end
			9062: begin bcd3<=9;bcd2<=0;bcd1<=6;bcd0<=2; end
			9063: begin bcd3<=9;bcd2<=0;bcd1<=6;bcd0<=3; end
			9064: begin bcd3<=9;bcd2<=0;bcd1<=6;bcd0<=4; end
			9065: begin bcd3<=9;bcd2<=0;bcd1<=6;bcd0<=5; end
			9066: begin bcd3<=9;bcd2<=0;bcd1<=6;bcd0<=6; end
			9067: begin bcd3<=9;bcd2<=0;bcd1<=6;bcd0<=7; end
			9068: begin bcd3<=9;bcd2<=0;bcd1<=6;bcd0<=8; end
			9069: begin bcd3<=9;bcd2<=0;bcd1<=6;bcd0<=9; end
			9070: begin bcd3<=9;bcd2<=0;bcd1<=7;bcd0<=0; end
			9071: begin bcd3<=9;bcd2<=0;bcd1<=7;bcd0<=1; end
			9072: begin bcd3<=9;bcd2<=0;bcd1<=7;bcd0<=2; end
			9073: begin bcd3<=9;bcd2<=0;bcd1<=7;bcd0<=3; end
			9074: begin bcd3<=9;bcd2<=0;bcd1<=7;bcd0<=4; end
			9075: begin bcd3<=9;bcd2<=0;bcd1<=7;bcd0<=5; end
			9076: begin bcd3<=9;bcd2<=0;bcd1<=7;bcd0<=6; end
			9077: begin bcd3<=9;bcd2<=0;bcd1<=7;bcd0<=7; end
			9078: begin bcd3<=9;bcd2<=0;bcd1<=7;bcd0<=8; end
			9079: begin bcd3<=9;bcd2<=0;bcd1<=7;bcd0<=9; end
			9080: begin bcd3<=9;bcd2<=0;bcd1<=8;bcd0<=0; end
			9081: begin bcd3<=9;bcd2<=0;bcd1<=8;bcd0<=1; end
			9082: begin bcd3<=9;bcd2<=0;bcd1<=8;bcd0<=2; end
			9083: begin bcd3<=9;bcd2<=0;bcd1<=8;bcd0<=3; end
			9084: begin bcd3<=9;bcd2<=0;bcd1<=8;bcd0<=4; end
			9085: begin bcd3<=9;bcd2<=0;bcd1<=8;bcd0<=5; end
			9086: begin bcd3<=9;bcd2<=0;bcd1<=8;bcd0<=6; end
			9087: begin bcd3<=9;bcd2<=0;bcd1<=8;bcd0<=7; end
			9088: begin bcd3<=9;bcd2<=0;bcd1<=8;bcd0<=8; end
			9089: begin bcd3<=9;bcd2<=0;bcd1<=8;bcd0<=9; end
			9090: begin bcd3<=9;bcd2<=0;bcd1<=9;bcd0<=0; end
			9091: begin bcd3<=9;bcd2<=0;bcd1<=9;bcd0<=1; end
			9092: begin bcd3<=9;bcd2<=0;bcd1<=9;bcd0<=2; end
			9093: begin bcd3<=9;bcd2<=0;bcd1<=9;bcd0<=3; end
			9094: begin bcd3<=9;bcd2<=0;bcd1<=9;bcd0<=4; end
			9095: begin bcd3<=9;bcd2<=0;bcd1<=9;bcd0<=5; end
			9096: begin bcd3<=9;bcd2<=0;bcd1<=9;bcd0<=6; end
			9097: begin bcd3<=9;bcd2<=0;bcd1<=9;bcd0<=7; end
			9098: begin bcd3<=9;bcd2<=0;bcd1<=9;bcd0<=8; end
			9099: begin bcd3<=9;bcd2<=0;bcd1<=9;bcd0<=9; end
			9100: begin bcd3<=9;bcd2<=1;bcd1<=0;bcd0<=0; end
			9101: begin bcd3<=9;bcd2<=1;bcd1<=0;bcd0<=1; end
			9102: begin bcd3<=9;bcd2<=1;bcd1<=0;bcd0<=2; end
			9103: begin bcd3<=9;bcd2<=1;bcd1<=0;bcd0<=3; end
			9104: begin bcd3<=9;bcd2<=1;bcd1<=0;bcd0<=4; end
			9105: begin bcd3<=9;bcd2<=1;bcd1<=0;bcd0<=5; end
			9106: begin bcd3<=9;bcd2<=1;bcd1<=0;bcd0<=6; end
			9107: begin bcd3<=9;bcd2<=1;bcd1<=0;bcd0<=7; end
			9108: begin bcd3<=9;bcd2<=1;bcd1<=0;bcd0<=8; end
			9109: begin bcd3<=9;bcd2<=1;bcd1<=0;bcd0<=9; end
			9110: begin bcd3<=9;bcd2<=1;bcd1<=1;bcd0<=0; end
			9111: begin bcd3<=9;bcd2<=1;bcd1<=1;bcd0<=1; end
			9112: begin bcd3<=9;bcd2<=1;bcd1<=1;bcd0<=2; end
			9113: begin bcd3<=9;bcd2<=1;bcd1<=1;bcd0<=3; end
			9114: begin bcd3<=9;bcd2<=1;bcd1<=1;bcd0<=4; end
			9115: begin bcd3<=9;bcd2<=1;bcd1<=1;bcd0<=5; end
			9116: begin bcd3<=9;bcd2<=1;bcd1<=1;bcd0<=6; end
			9117: begin bcd3<=9;bcd2<=1;bcd1<=1;bcd0<=7; end
			9118: begin bcd3<=9;bcd2<=1;bcd1<=1;bcd0<=8; end
			9119: begin bcd3<=9;bcd2<=1;bcd1<=1;bcd0<=9; end
			9120: begin bcd3<=9;bcd2<=1;bcd1<=2;bcd0<=0; end
			9121: begin bcd3<=9;bcd2<=1;bcd1<=2;bcd0<=1; end
			9122: begin bcd3<=9;bcd2<=1;bcd1<=2;bcd0<=2; end
			9123: begin bcd3<=9;bcd2<=1;bcd1<=2;bcd0<=3; end
			9124: begin bcd3<=9;bcd2<=1;bcd1<=2;bcd0<=4; end
			9125: begin bcd3<=9;bcd2<=1;bcd1<=2;bcd0<=5; end
			9126: begin bcd3<=9;bcd2<=1;bcd1<=2;bcd0<=6; end
			9127: begin bcd3<=9;bcd2<=1;bcd1<=2;bcd0<=7; end
			9128: begin bcd3<=9;bcd2<=1;bcd1<=2;bcd0<=8; end
			9129: begin bcd3<=9;bcd2<=1;bcd1<=2;bcd0<=9; end
			9130: begin bcd3<=9;bcd2<=1;bcd1<=3;bcd0<=0; end
			9131: begin bcd3<=9;bcd2<=1;bcd1<=3;bcd0<=1; end
			9132: begin bcd3<=9;bcd2<=1;bcd1<=3;bcd0<=2; end
			9133: begin bcd3<=9;bcd2<=1;bcd1<=3;bcd0<=3; end
			9134: begin bcd3<=9;bcd2<=1;bcd1<=3;bcd0<=4; end
			9135: begin bcd3<=9;bcd2<=1;bcd1<=3;bcd0<=5; end
			9136: begin bcd3<=9;bcd2<=1;bcd1<=3;bcd0<=6; end
			9137: begin bcd3<=9;bcd2<=1;bcd1<=3;bcd0<=7; end
			9138: begin bcd3<=9;bcd2<=1;bcd1<=3;bcd0<=8; end
			9139: begin bcd3<=9;bcd2<=1;bcd1<=3;bcd0<=9; end
			9140: begin bcd3<=9;bcd2<=1;bcd1<=4;bcd0<=0; end
			9141: begin bcd3<=9;bcd2<=1;bcd1<=4;bcd0<=1; end
			9142: begin bcd3<=9;bcd2<=1;bcd1<=4;bcd0<=2; end
			9143: begin bcd3<=9;bcd2<=1;bcd1<=4;bcd0<=3; end
			9144: begin bcd3<=9;bcd2<=1;bcd1<=4;bcd0<=4; end
			9145: begin bcd3<=9;bcd2<=1;bcd1<=4;bcd0<=5; end
			9146: begin bcd3<=9;bcd2<=1;bcd1<=4;bcd0<=6; end
			9147: begin bcd3<=9;bcd2<=1;bcd1<=4;bcd0<=7; end
			9148: begin bcd3<=9;bcd2<=1;bcd1<=4;bcd0<=8; end
			9149: begin bcd3<=9;bcd2<=1;bcd1<=4;bcd0<=9; end
			9150: begin bcd3<=9;bcd2<=1;bcd1<=5;bcd0<=0; end
			9151: begin bcd3<=9;bcd2<=1;bcd1<=5;bcd0<=1; end
			9152: begin bcd3<=9;bcd2<=1;bcd1<=5;bcd0<=2; end
			9153: begin bcd3<=9;bcd2<=1;bcd1<=5;bcd0<=3; end
			9154: begin bcd3<=9;bcd2<=1;bcd1<=5;bcd0<=4; end
			9155: begin bcd3<=9;bcd2<=1;bcd1<=5;bcd0<=5; end
			9156: begin bcd3<=9;bcd2<=1;bcd1<=5;bcd0<=6; end
			9157: begin bcd3<=9;bcd2<=1;bcd1<=5;bcd0<=7; end
			9158: begin bcd3<=9;bcd2<=1;bcd1<=5;bcd0<=8; end
			9159: begin bcd3<=9;bcd2<=1;bcd1<=5;bcd0<=9; end
			9160: begin bcd3<=9;bcd2<=1;bcd1<=6;bcd0<=0; end
			9161: begin bcd3<=9;bcd2<=1;bcd1<=6;bcd0<=1; end
			9162: begin bcd3<=9;bcd2<=1;bcd1<=6;bcd0<=2; end
			9163: begin bcd3<=9;bcd2<=1;bcd1<=6;bcd0<=3; end
			9164: begin bcd3<=9;bcd2<=1;bcd1<=6;bcd0<=4; end
			9165: begin bcd3<=9;bcd2<=1;bcd1<=6;bcd0<=5; end
			9166: begin bcd3<=9;bcd2<=1;bcd1<=6;bcd0<=6; end
			9167: begin bcd3<=9;bcd2<=1;bcd1<=6;bcd0<=7; end
			9168: begin bcd3<=9;bcd2<=1;bcd1<=6;bcd0<=8; end
			9169: begin bcd3<=9;bcd2<=1;bcd1<=6;bcd0<=9; end
			9170: begin bcd3<=9;bcd2<=1;bcd1<=7;bcd0<=0; end
			9171: begin bcd3<=9;bcd2<=1;bcd1<=7;bcd0<=1; end
			9172: begin bcd3<=9;bcd2<=1;bcd1<=7;bcd0<=2; end
			9173: begin bcd3<=9;bcd2<=1;bcd1<=7;bcd0<=3; end
			9174: begin bcd3<=9;bcd2<=1;bcd1<=7;bcd0<=4; end
			9175: begin bcd3<=9;bcd2<=1;bcd1<=7;bcd0<=5; end
			9176: begin bcd3<=9;bcd2<=1;bcd1<=7;bcd0<=6; end
			9177: begin bcd3<=9;bcd2<=1;bcd1<=7;bcd0<=7; end
			9178: begin bcd3<=9;bcd2<=1;bcd1<=7;bcd0<=8; end
			9179: begin bcd3<=9;bcd2<=1;bcd1<=7;bcd0<=9; end
			9180: begin bcd3<=9;bcd2<=1;bcd1<=8;bcd0<=0; end
			9181: begin bcd3<=9;bcd2<=1;bcd1<=8;bcd0<=1; end
			9182: begin bcd3<=9;bcd2<=1;bcd1<=8;bcd0<=2; end
			9183: begin bcd3<=9;bcd2<=1;bcd1<=8;bcd0<=3; end
			9184: begin bcd3<=9;bcd2<=1;bcd1<=8;bcd0<=4; end
			9185: begin bcd3<=9;bcd2<=1;bcd1<=8;bcd0<=5; end
			9186: begin bcd3<=9;bcd2<=1;bcd1<=8;bcd0<=6; end
			9187: begin bcd3<=9;bcd2<=1;bcd1<=8;bcd0<=7; end
			9188: begin bcd3<=9;bcd2<=1;bcd1<=8;bcd0<=8; end
			9189: begin bcd3<=9;bcd2<=1;bcd1<=8;bcd0<=9; end
			9190: begin bcd3<=9;bcd2<=1;bcd1<=9;bcd0<=0; end
			9191: begin bcd3<=9;bcd2<=1;bcd1<=9;bcd0<=1; end
			9192: begin bcd3<=9;bcd2<=1;bcd1<=9;bcd0<=2; end
			9193: begin bcd3<=9;bcd2<=1;bcd1<=9;bcd0<=3; end
			9194: begin bcd3<=9;bcd2<=1;bcd1<=9;bcd0<=4; end
			9195: begin bcd3<=9;bcd2<=1;bcd1<=9;bcd0<=5; end
			9196: begin bcd3<=9;bcd2<=1;bcd1<=9;bcd0<=6; end
			9197: begin bcd3<=9;bcd2<=1;bcd1<=9;bcd0<=7; end
			9198: begin bcd3<=9;bcd2<=1;bcd1<=9;bcd0<=8; end
			9199: begin bcd3<=9;bcd2<=1;bcd1<=9;bcd0<=9; end
			9200: begin bcd3<=9;bcd2<=2;bcd1<=0;bcd0<=0; end
			9201: begin bcd3<=9;bcd2<=2;bcd1<=0;bcd0<=1; end
			9202: begin bcd3<=9;bcd2<=2;bcd1<=0;bcd0<=2; end
			9203: begin bcd3<=9;bcd2<=2;bcd1<=0;bcd0<=3; end
			9204: begin bcd3<=9;bcd2<=2;bcd1<=0;bcd0<=4; end
			9205: begin bcd3<=9;bcd2<=2;bcd1<=0;bcd0<=5; end
			9206: begin bcd3<=9;bcd2<=2;bcd1<=0;bcd0<=6; end
			9207: begin bcd3<=9;bcd2<=2;bcd1<=0;bcd0<=7; end
			9208: begin bcd3<=9;bcd2<=2;bcd1<=0;bcd0<=8; end
			9209: begin bcd3<=9;bcd2<=2;bcd1<=0;bcd0<=9; end
			9210: begin bcd3<=9;bcd2<=2;bcd1<=1;bcd0<=0; end
			9211: begin bcd3<=9;bcd2<=2;bcd1<=1;bcd0<=1; end
			9212: begin bcd3<=9;bcd2<=2;bcd1<=1;bcd0<=2; end
			9213: begin bcd3<=9;bcd2<=2;bcd1<=1;bcd0<=3; end
			9214: begin bcd3<=9;bcd2<=2;bcd1<=1;bcd0<=4; end
			9215: begin bcd3<=9;bcd2<=2;bcd1<=1;bcd0<=5; end
			9216: begin bcd3<=9;bcd2<=2;bcd1<=1;bcd0<=6; end
			9217: begin bcd3<=9;bcd2<=2;bcd1<=1;bcd0<=7; end
			9218: begin bcd3<=9;bcd2<=2;bcd1<=1;bcd0<=8; end
			9219: begin bcd3<=9;bcd2<=2;bcd1<=1;bcd0<=9; end
			9220: begin bcd3<=9;bcd2<=2;bcd1<=2;bcd0<=0; end
			9221: begin bcd3<=9;bcd2<=2;bcd1<=2;bcd0<=1; end
			9222: begin bcd3<=9;bcd2<=2;bcd1<=2;bcd0<=2; end
			9223: begin bcd3<=9;bcd2<=2;bcd1<=2;bcd0<=3; end
			9224: begin bcd3<=9;bcd2<=2;bcd1<=2;bcd0<=4; end
			9225: begin bcd3<=9;bcd2<=2;bcd1<=2;bcd0<=5; end
			9226: begin bcd3<=9;bcd2<=2;bcd1<=2;bcd0<=6; end
			9227: begin bcd3<=9;bcd2<=2;bcd1<=2;bcd0<=7; end
			9228: begin bcd3<=9;bcd2<=2;bcd1<=2;bcd0<=8; end
			9229: begin bcd3<=9;bcd2<=2;bcd1<=2;bcd0<=9; end
			9230: begin bcd3<=9;bcd2<=2;bcd1<=3;bcd0<=0; end
			9231: begin bcd3<=9;bcd2<=2;bcd1<=3;bcd0<=1; end
			9232: begin bcd3<=9;bcd2<=2;bcd1<=3;bcd0<=2; end
			9233: begin bcd3<=9;bcd2<=2;bcd1<=3;bcd0<=3; end
			9234: begin bcd3<=9;bcd2<=2;bcd1<=3;bcd0<=4; end
			9235: begin bcd3<=9;bcd2<=2;bcd1<=3;bcd0<=5; end
			9236: begin bcd3<=9;bcd2<=2;bcd1<=3;bcd0<=6; end
			9237: begin bcd3<=9;bcd2<=2;bcd1<=3;bcd0<=7; end
			9238: begin bcd3<=9;bcd2<=2;bcd1<=3;bcd0<=8; end
			9239: begin bcd3<=9;bcd2<=2;bcd1<=3;bcd0<=9; end
			9240: begin bcd3<=9;bcd2<=2;bcd1<=4;bcd0<=0; end
			9241: begin bcd3<=9;bcd2<=2;bcd1<=4;bcd0<=1; end
			9242: begin bcd3<=9;bcd2<=2;bcd1<=4;bcd0<=2; end
			9243: begin bcd3<=9;bcd2<=2;bcd1<=4;bcd0<=3; end
			9244: begin bcd3<=9;bcd2<=2;bcd1<=4;bcd0<=4; end
			9245: begin bcd3<=9;bcd2<=2;bcd1<=4;bcd0<=5; end
			9246: begin bcd3<=9;bcd2<=2;bcd1<=4;bcd0<=6; end
			9247: begin bcd3<=9;bcd2<=2;bcd1<=4;bcd0<=7; end
			9248: begin bcd3<=9;bcd2<=2;bcd1<=4;bcd0<=8; end
			9249: begin bcd3<=9;bcd2<=2;bcd1<=4;bcd0<=9; end
			9250: begin bcd3<=9;bcd2<=2;bcd1<=5;bcd0<=0; end
			9251: begin bcd3<=9;bcd2<=2;bcd1<=5;bcd0<=1; end
			9252: begin bcd3<=9;bcd2<=2;bcd1<=5;bcd0<=2; end
			9253: begin bcd3<=9;bcd2<=2;bcd1<=5;bcd0<=3; end
			9254: begin bcd3<=9;bcd2<=2;bcd1<=5;bcd0<=4; end
			9255: begin bcd3<=9;bcd2<=2;bcd1<=5;bcd0<=5; end
			9256: begin bcd3<=9;bcd2<=2;bcd1<=5;bcd0<=6; end
			9257: begin bcd3<=9;bcd2<=2;bcd1<=5;bcd0<=7; end
			9258: begin bcd3<=9;bcd2<=2;bcd1<=5;bcd0<=8; end
			9259: begin bcd3<=9;bcd2<=2;bcd1<=5;bcd0<=9; end
			9260: begin bcd3<=9;bcd2<=2;bcd1<=6;bcd0<=0; end
			9261: begin bcd3<=9;bcd2<=2;bcd1<=6;bcd0<=1; end
			9262: begin bcd3<=9;bcd2<=2;bcd1<=6;bcd0<=2; end
			9263: begin bcd3<=9;bcd2<=2;bcd1<=6;bcd0<=3; end
			9264: begin bcd3<=9;bcd2<=2;bcd1<=6;bcd0<=4; end
			9265: begin bcd3<=9;bcd2<=2;bcd1<=6;bcd0<=5; end
			9266: begin bcd3<=9;bcd2<=2;bcd1<=6;bcd0<=6; end
			9267: begin bcd3<=9;bcd2<=2;bcd1<=6;bcd0<=7; end
			9268: begin bcd3<=9;bcd2<=2;bcd1<=6;bcd0<=8; end
			9269: begin bcd3<=9;bcd2<=2;bcd1<=6;bcd0<=9; end
			9270: begin bcd3<=9;bcd2<=2;bcd1<=7;bcd0<=0; end
			9271: begin bcd3<=9;bcd2<=2;bcd1<=7;bcd0<=1; end
			9272: begin bcd3<=9;bcd2<=2;bcd1<=7;bcd0<=2; end
			9273: begin bcd3<=9;bcd2<=2;bcd1<=7;bcd0<=3; end
			9274: begin bcd3<=9;bcd2<=2;bcd1<=7;bcd0<=4; end
			9275: begin bcd3<=9;bcd2<=2;bcd1<=7;bcd0<=5; end
			9276: begin bcd3<=9;bcd2<=2;bcd1<=7;bcd0<=6; end
			9277: begin bcd3<=9;bcd2<=2;bcd1<=7;bcd0<=7; end
			9278: begin bcd3<=9;bcd2<=2;bcd1<=7;bcd0<=8; end
			9279: begin bcd3<=9;bcd2<=2;bcd1<=7;bcd0<=9; end
			9280: begin bcd3<=9;bcd2<=2;bcd1<=8;bcd0<=0; end
			9281: begin bcd3<=9;bcd2<=2;bcd1<=8;bcd0<=1; end
			9282: begin bcd3<=9;bcd2<=2;bcd1<=8;bcd0<=2; end
			9283: begin bcd3<=9;bcd2<=2;bcd1<=8;bcd0<=3; end
			9284: begin bcd3<=9;bcd2<=2;bcd1<=8;bcd0<=4; end
			9285: begin bcd3<=9;bcd2<=2;bcd1<=8;bcd0<=5; end
			9286: begin bcd3<=9;bcd2<=2;bcd1<=8;bcd0<=6; end
			9287: begin bcd3<=9;bcd2<=2;bcd1<=8;bcd0<=7; end
			9288: begin bcd3<=9;bcd2<=2;bcd1<=8;bcd0<=8; end
			9289: begin bcd3<=9;bcd2<=2;bcd1<=8;bcd0<=9; end
			9290: begin bcd3<=9;bcd2<=2;bcd1<=9;bcd0<=0; end
			9291: begin bcd3<=9;bcd2<=2;bcd1<=9;bcd0<=1; end
			9292: begin bcd3<=9;bcd2<=2;bcd1<=9;bcd0<=2; end
			9293: begin bcd3<=9;bcd2<=2;bcd1<=9;bcd0<=3; end
			9294: begin bcd3<=9;bcd2<=2;bcd1<=9;bcd0<=4; end
			9295: begin bcd3<=9;bcd2<=2;bcd1<=9;bcd0<=5; end
			9296: begin bcd3<=9;bcd2<=2;bcd1<=9;bcd0<=6; end
			9297: begin bcd3<=9;bcd2<=2;bcd1<=9;bcd0<=7; end
			9298: begin bcd3<=9;bcd2<=2;bcd1<=9;bcd0<=8; end
			9299: begin bcd3<=9;bcd2<=2;bcd1<=9;bcd0<=9; end
			9300: begin bcd3<=9;bcd2<=3;bcd1<=0;bcd0<=0; end
			9301: begin bcd3<=9;bcd2<=3;bcd1<=0;bcd0<=1; end
			9302: begin bcd3<=9;bcd2<=3;bcd1<=0;bcd0<=2; end
			9303: begin bcd3<=9;bcd2<=3;bcd1<=0;bcd0<=3; end
			9304: begin bcd3<=9;bcd2<=3;bcd1<=0;bcd0<=4; end
			9305: begin bcd3<=9;bcd2<=3;bcd1<=0;bcd0<=5; end
			9306: begin bcd3<=9;bcd2<=3;bcd1<=0;bcd0<=6; end
			9307: begin bcd3<=9;bcd2<=3;bcd1<=0;bcd0<=7; end
			9308: begin bcd3<=9;bcd2<=3;bcd1<=0;bcd0<=8; end
			9309: begin bcd3<=9;bcd2<=3;bcd1<=0;bcd0<=9; end
			9310: begin bcd3<=9;bcd2<=3;bcd1<=1;bcd0<=0; end
			9311: begin bcd3<=9;bcd2<=3;bcd1<=1;bcd0<=1; end
			9312: begin bcd3<=9;bcd2<=3;bcd1<=1;bcd0<=2; end
			9313: begin bcd3<=9;bcd2<=3;bcd1<=1;bcd0<=3; end
			9314: begin bcd3<=9;bcd2<=3;bcd1<=1;bcd0<=4; end
			9315: begin bcd3<=9;bcd2<=3;bcd1<=1;bcd0<=5; end
			9316: begin bcd3<=9;bcd2<=3;bcd1<=1;bcd0<=6; end
			9317: begin bcd3<=9;bcd2<=3;bcd1<=1;bcd0<=7; end
			9318: begin bcd3<=9;bcd2<=3;bcd1<=1;bcd0<=8; end
			9319: begin bcd3<=9;bcd2<=3;bcd1<=1;bcd0<=9; end
			9320: begin bcd3<=9;bcd2<=3;bcd1<=2;bcd0<=0; end
			9321: begin bcd3<=9;bcd2<=3;bcd1<=2;bcd0<=1; end
			9322: begin bcd3<=9;bcd2<=3;bcd1<=2;bcd0<=2; end
			9323: begin bcd3<=9;bcd2<=3;bcd1<=2;bcd0<=3; end
			9324: begin bcd3<=9;bcd2<=3;bcd1<=2;bcd0<=4; end
			9325: begin bcd3<=9;bcd2<=3;bcd1<=2;bcd0<=5; end
			9326: begin bcd3<=9;bcd2<=3;bcd1<=2;bcd0<=6; end
			9327: begin bcd3<=9;bcd2<=3;bcd1<=2;bcd0<=7; end
			9328: begin bcd3<=9;bcd2<=3;bcd1<=2;bcd0<=8; end
			9329: begin bcd3<=9;bcd2<=3;bcd1<=2;bcd0<=9; end
			9330: begin bcd3<=9;bcd2<=3;bcd1<=3;bcd0<=0; end
			9331: begin bcd3<=9;bcd2<=3;bcd1<=3;bcd0<=1; end
			9332: begin bcd3<=9;bcd2<=3;bcd1<=3;bcd0<=2; end
			9333: begin bcd3<=9;bcd2<=3;bcd1<=3;bcd0<=3; end
			9334: begin bcd3<=9;bcd2<=3;bcd1<=3;bcd0<=4; end
			9335: begin bcd3<=9;bcd2<=3;bcd1<=3;bcd0<=5; end
			9336: begin bcd3<=9;bcd2<=3;bcd1<=3;bcd0<=6; end
			9337: begin bcd3<=9;bcd2<=3;bcd1<=3;bcd0<=7; end
			9338: begin bcd3<=9;bcd2<=3;bcd1<=3;bcd0<=8; end
			9339: begin bcd3<=9;bcd2<=3;bcd1<=3;bcd0<=9; end
			9340: begin bcd3<=9;bcd2<=3;bcd1<=4;bcd0<=0; end
			9341: begin bcd3<=9;bcd2<=3;bcd1<=4;bcd0<=1; end
			9342: begin bcd3<=9;bcd2<=3;bcd1<=4;bcd0<=2; end
			9343: begin bcd3<=9;bcd2<=3;bcd1<=4;bcd0<=3; end
			9344: begin bcd3<=9;bcd2<=3;bcd1<=4;bcd0<=4; end
			9345: begin bcd3<=9;bcd2<=3;bcd1<=4;bcd0<=5; end
			9346: begin bcd3<=9;bcd2<=3;bcd1<=4;bcd0<=6; end
			9347: begin bcd3<=9;bcd2<=3;bcd1<=4;bcd0<=7; end
			9348: begin bcd3<=9;bcd2<=3;bcd1<=4;bcd0<=8; end
			9349: begin bcd3<=9;bcd2<=3;bcd1<=4;bcd0<=9; end
			9350: begin bcd3<=9;bcd2<=3;bcd1<=5;bcd0<=0; end
			9351: begin bcd3<=9;bcd2<=3;bcd1<=5;bcd0<=1; end
			9352: begin bcd3<=9;bcd2<=3;bcd1<=5;bcd0<=2; end
			9353: begin bcd3<=9;bcd2<=3;bcd1<=5;bcd0<=3; end
			9354: begin bcd3<=9;bcd2<=3;bcd1<=5;bcd0<=4; end
			9355: begin bcd3<=9;bcd2<=3;bcd1<=5;bcd0<=5; end
			9356: begin bcd3<=9;bcd2<=3;bcd1<=5;bcd0<=6; end
			9357: begin bcd3<=9;bcd2<=3;bcd1<=5;bcd0<=7; end
			9358: begin bcd3<=9;bcd2<=3;bcd1<=5;bcd0<=8; end
			9359: begin bcd3<=9;bcd2<=3;bcd1<=5;bcd0<=9; end
			9360: begin bcd3<=9;bcd2<=3;bcd1<=6;bcd0<=0; end
			9361: begin bcd3<=9;bcd2<=3;bcd1<=6;bcd0<=1; end
			9362: begin bcd3<=9;bcd2<=3;bcd1<=6;bcd0<=2; end
			9363: begin bcd3<=9;bcd2<=3;bcd1<=6;bcd0<=3; end
			9364: begin bcd3<=9;bcd2<=3;bcd1<=6;bcd0<=4; end
			9365: begin bcd3<=9;bcd2<=3;bcd1<=6;bcd0<=5; end
			9366: begin bcd3<=9;bcd2<=3;bcd1<=6;bcd0<=6; end
			9367: begin bcd3<=9;bcd2<=3;bcd1<=6;bcd0<=7; end
			9368: begin bcd3<=9;bcd2<=3;bcd1<=6;bcd0<=8; end
			9369: begin bcd3<=9;bcd2<=3;bcd1<=6;bcd0<=9; end
			9370: begin bcd3<=9;bcd2<=3;bcd1<=7;bcd0<=0; end
			9371: begin bcd3<=9;bcd2<=3;bcd1<=7;bcd0<=1; end
			9372: begin bcd3<=9;bcd2<=3;bcd1<=7;bcd0<=2; end
			9373: begin bcd3<=9;bcd2<=3;bcd1<=7;bcd0<=3; end
			9374: begin bcd3<=9;bcd2<=3;bcd1<=7;bcd0<=4; end
			9375: begin bcd3<=9;bcd2<=3;bcd1<=7;bcd0<=5; end
			9376: begin bcd3<=9;bcd2<=3;bcd1<=7;bcd0<=6; end
			9377: begin bcd3<=9;bcd2<=3;bcd1<=7;bcd0<=7; end
			9378: begin bcd3<=9;bcd2<=3;bcd1<=7;bcd0<=8; end
			9379: begin bcd3<=9;bcd2<=3;bcd1<=7;bcd0<=9; end
			9380: begin bcd3<=9;bcd2<=3;bcd1<=8;bcd0<=0; end
			9381: begin bcd3<=9;bcd2<=3;bcd1<=8;bcd0<=1; end
			9382: begin bcd3<=9;bcd2<=3;bcd1<=8;bcd0<=2; end
			9383: begin bcd3<=9;bcd2<=3;bcd1<=8;bcd0<=3; end
			9384: begin bcd3<=9;bcd2<=3;bcd1<=8;bcd0<=4; end
			9385: begin bcd3<=9;bcd2<=3;bcd1<=8;bcd0<=5; end
			9386: begin bcd3<=9;bcd2<=3;bcd1<=8;bcd0<=6; end
			9387: begin bcd3<=9;bcd2<=3;bcd1<=8;bcd0<=7; end
			9388: begin bcd3<=9;bcd2<=3;bcd1<=8;bcd0<=8; end
			9389: begin bcd3<=9;bcd2<=3;bcd1<=8;bcd0<=9; end
			9390: begin bcd3<=9;bcd2<=3;bcd1<=9;bcd0<=0; end
			9391: begin bcd3<=9;bcd2<=3;bcd1<=9;bcd0<=1; end
			9392: begin bcd3<=9;bcd2<=3;bcd1<=9;bcd0<=2; end
			9393: begin bcd3<=9;bcd2<=3;bcd1<=9;bcd0<=3; end
			9394: begin bcd3<=9;bcd2<=3;bcd1<=9;bcd0<=4; end
			9395: begin bcd3<=9;bcd2<=3;bcd1<=9;bcd0<=5; end
			9396: begin bcd3<=9;bcd2<=3;bcd1<=9;bcd0<=6; end
			9397: begin bcd3<=9;bcd2<=3;bcd1<=9;bcd0<=7; end
			9398: begin bcd3<=9;bcd2<=3;bcd1<=9;bcd0<=8; end
			9399: begin bcd3<=9;bcd2<=3;bcd1<=9;bcd0<=9; end
			9400: begin bcd3<=9;bcd2<=4;bcd1<=0;bcd0<=0; end
			9401: begin bcd3<=9;bcd2<=4;bcd1<=0;bcd0<=1; end
			9402: begin bcd3<=9;bcd2<=4;bcd1<=0;bcd0<=2; end
			9403: begin bcd3<=9;bcd2<=4;bcd1<=0;bcd0<=3; end
			9404: begin bcd3<=9;bcd2<=4;bcd1<=0;bcd0<=4; end
			9405: begin bcd3<=9;bcd2<=4;bcd1<=0;bcd0<=5; end
			9406: begin bcd3<=9;bcd2<=4;bcd1<=0;bcd0<=6; end
			9407: begin bcd3<=9;bcd2<=4;bcd1<=0;bcd0<=7; end
			9408: begin bcd3<=9;bcd2<=4;bcd1<=0;bcd0<=8; end
			9409: begin bcd3<=9;bcd2<=4;bcd1<=0;bcd0<=9; end
			9410: begin bcd3<=9;bcd2<=4;bcd1<=1;bcd0<=0; end
			9411: begin bcd3<=9;bcd2<=4;bcd1<=1;bcd0<=1; end
			9412: begin bcd3<=9;bcd2<=4;bcd1<=1;bcd0<=2; end
			9413: begin bcd3<=9;bcd2<=4;bcd1<=1;bcd0<=3; end
			9414: begin bcd3<=9;bcd2<=4;bcd1<=1;bcd0<=4; end
			9415: begin bcd3<=9;bcd2<=4;bcd1<=1;bcd0<=5; end
			9416: begin bcd3<=9;bcd2<=4;bcd1<=1;bcd0<=6; end
			9417: begin bcd3<=9;bcd2<=4;bcd1<=1;bcd0<=7; end
			9418: begin bcd3<=9;bcd2<=4;bcd1<=1;bcd0<=8; end
			9419: begin bcd3<=9;bcd2<=4;bcd1<=1;bcd0<=9; end
			9420: begin bcd3<=9;bcd2<=4;bcd1<=2;bcd0<=0; end
			9421: begin bcd3<=9;bcd2<=4;bcd1<=2;bcd0<=1; end
			9422: begin bcd3<=9;bcd2<=4;bcd1<=2;bcd0<=2; end
			9423: begin bcd3<=9;bcd2<=4;bcd1<=2;bcd0<=3; end
			9424: begin bcd3<=9;bcd2<=4;bcd1<=2;bcd0<=4; end
			9425: begin bcd3<=9;bcd2<=4;bcd1<=2;bcd0<=5; end
			9426: begin bcd3<=9;bcd2<=4;bcd1<=2;bcd0<=6; end
			9427: begin bcd3<=9;bcd2<=4;bcd1<=2;bcd0<=7; end
			9428: begin bcd3<=9;bcd2<=4;bcd1<=2;bcd0<=8; end
			9429: begin bcd3<=9;bcd2<=4;bcd1<=2;bcd0<=9; end
			9430: begin bcd3<=9;bcd2<=4;bcd1<=3;bcd0<=0; end
			9431: begin bcd3<=9;bcd2<=4;bcd1<=3;bcd0<=1; end
			9432: begin bcd3<=9;bcd2<=4;bcd1<=3;bcd0<=2; end
			9433: begin bcd3<=9;bcd2<=4;bcd1<=3;bcd0<=3; end
			9434: begin bcd3<=9;bcd2<=4;bcd1<=3;bcd0<=4; end
			9435: begin bcd3<=9;bcd2<=4;bcd1<=3;bcd0<=5; end
			9436: begin bcd3<=9;bcd2<=4;bcd1<=3;bcd0<=6; end
			9437: begin bcd3<=9;bcd2<=4;bcd1<=3;bcd0<=7; end
			9438: begin bcd3<=9;bcd2<=4;bcd1<=3;bcd0<=8; end
			9439: begin bcd3<=9;bcd2<=4;bcd1<=3;bcd0<=9; end
			9440: begin bcd3<=9;bcd2<=4;bcd1<=4;bcd0<=0; end
			9441: begin bcd3<=9;bcd2<=4;bcd1<=4;bcd0<=1; end
			9442: begin bcd3<=9;bcd2<=4;bcd1<=4;bcd0<=2; end
			9443: begin bcd3<=9;bcd2<=4;bcd1<=4;bcd0<=3; end
			9444: begin bcd3<=9;bcd2<=4;bcd1<=4;bcd0<=4; end
			9445: begin bcd3<=9;bcd2<=4;bcd1<=4;bcd0<=5; end
			9446: begin bcd3<=9;bcd2<=4;bcd1<=4;bcd0<=6; end
			9447: begin bcd3<=9;bcd2<=4;bcd1<=4;bcd0<=7; end
			9448: begin bcd3<=9;bcd2<=4;bcd1<=4;bcd0<=8; end
			9449: begin bcd3<=9;bcd2<=4;bcd1<=4;bcd0<=9; end
			9450: begin bcd3<=9;bcd2<=4;bcd1<=5;bcd0<=0; end
			9451: begin bcd3<=9;bcd2<=4;bcd1<=5;bcd0<=1; end
			9452: begin bcd3<=9;bcd2<=4;bcd1<=5;bcd0<=2; end
			9453: begin bcd3<=9;bcd2<=4;bcd1<=5;bcd0<=3; end
			9454: begin bcd3<=9;bcd2<=4;bcd1<=5;bcd0<=4; end
			9455: begin bcd3<=9;bcd2<=4;bcd1<=5;bcd0<=5; end
			9456: begin bcd3<=9;bcd2<=4;bcd1<=5;bcd0<=6; end
			9457: begin bcd3<=9;bcd2<=4;bcd1<=5;bcd0<=7; end
			9458: begin bcd3<=9;bcd2<=4;bcd1<=5;bcd0<=8; end
			9459: begin bcd3<=9;bcd2<=4;bcd1<=5;bcd0<=9; end
			9460: begin bcd3<=9;bcd2<=4;bcd1<=6;bcd0<=0; end
			9461: begin bcd3<=9;bcd2<=4;bcd1<=6;bcd0<=1; end
			9462: begin bcd3<=9;bcd2<=4;bcd1<=6;bcd0<=2; end
			9463: begin bcd3<=9;bcd2<=4;bcd1<=6;bcd0<=3; end
			9464: begin bcd3<=9;bcd2<=4;bcd1<=6;bcd0<=4; end
			9465: begin bcd3<=9;bcd2<=4;bcd1<=6;bcd0<=5; end
			9466: begin bcd3<=9;bcd2<=4;bcd1<=6;bcd0<=6; end
			9467: begin bcd3<=9;bcd2<=4;bcd1<=6;bcd0<=7; end
			9468: begin bcd3<=9;bcd2<=4;bcd1<=6;bcd0<=8; end
			9469: begin bcd3<=9;bcd2<=4;bcd1<=6;bcd0<=9; end
			9470: begin bcd3<=9;bcd2<=4;bcd1<=7;bcd0<=0; end
			9471: begin bcd3<=9;bcd2<=4;bcd1<=7;bcd0<=1; end
			9472: begin bcd3<=9;bcd2<=4;bcd1<=7;bcd0<=2; end
			9473: begin bcd3<=9;bcd2<=4;bcd1<=7;bcd0<=3; end
			9474: begin bcd3<=9;bcd2<=4;bcd1<=7;bcd0<=4; end
			9475: begin bcd3<=9;bcd2<=4;bcd1<=7;bcd0<=5; end
			9476: begin bcd3<=9;bcd2<=4;bcd1<=7;bcd0<=6; end
			9477: begin bcd3<=9;bcd2<=4;bcd1<=7;bcd0<=7; end
			9478: begin bcd3<=9;bcd2<=4;bcd1<=7;bcd0<=8; end
			9479: begin bcd3<=9;bcd2<=4;bcd1<=7;bcd0<=9; end
			9480: begin bcd3<=9;bcd2<=4;bcd1<=8;bcd0<=0; end
			9481: begin bcd3<=9;bcd2<=4;bcd1<=8;bcd0<=1; end
			9482: begin bcd3<=9;bcd2<=4;bcd1<=8;bcd0<=2; end
			9483: begin bcd3<=9;bcd2<=4;bcd1<=8;bcd0<=3; end
			9484: begin bcd3<=9;bcd2<=4;bcd1<=8;bcd0<=4; end
			9485: begin bcd3<=9;bcd2<=4;bcd1<=8;bcd0<=5; end
			9486: begin bcd3<=9;bcd2<=4;bcd1<=8;bcd0<=6; end
			9487: begin bcd3<=9;bcd2<=4;bcd1<=8;bcd0<=7; end
			9488: begin bcd3<=9;bcd2<=4;bcd1<=8;bcd0<=8; end
			9489: begin bcd3<=9;bcd2<=4;bcd1<=8;bcd0<=9; end
			9490: begin bcd3<=9;bcd2<=4;bcd1<=9;bcd0<=0; end
			9491: begin bcd3<=9;bcd2<=4;bcd1<=9;bcd0<=1; end
			9492: begin bcd3<=9;bcd2<=4;bcd1<=9;bcd0<=2; end
			9493: begin bcd3<=9;bcd2<=4;bcd1<=9;bcd0<=3; end
			9494: begin bcd3<=9;bcd2<=4;bcd1<=9;bcd0<=4; end
			9495: begin bcd3<=9;bcd2<=4;bcd1<=9;bcd0<=5; end
			9496: begin bcd3<=9;bcd2<=4;bcd1<=9;bcd0<=6; end
			9497: begin bcd3<=9;bcd2<=4;bcd1<=9;bcd0<=7; end
			9498: begin bcd3<=9;bcd2<=4;bcd1<=9;bcd0<=8; end
			9499: begin bcd3<=9;bcd2<=4;bcd1<=9;bcd0<=9; end
			9500: begin bcd3<=9;bcd2<=5;bcd1<=0;bcd0<=0; end
			9501: begin bcd3<=9;bcd2<=5;bcd1<=0;bcd0<=1; end
			9502: begin bcd3<=9;bcd2<=5;bcd1<=0;bcd0<=2; end
			9503: begin bcd3<=9;bcd2<=5;bcd1<=0;bcd0<=3; end
			9504: begin bcd3<=9;bcd2<=5;bcd1<=0;bcd0<=4; end
			9505: begin bcd3<=9;bcd2<=5;bcd1<=0;bcd0<=5; end
			9506: begin bcd3<=9;bcd2<=5;bcd1<=0;bcd0<=6; end
			9507: begin bcd3<=9;bcd2<=5;bcd1<=0;bcd0<=7; end
			9508: begin bcd3<=9;bcd2<=5;bcd1<=0;bcd0<=8; end
			9509: begin bcd3<=9;bcd2<=5;bcd1<=0;bcd0<=9; end
			9510: begin bcd3<=9;bcd2<=5;bcd1<=1;bcd0<=0; end
			9511: begin bcd3<=9;bcd2<=5;bcd1<=1;bcd0<=1; end
			9512: begin bcd3<=9;bcd2<=5;bcd1<=1;bcd0<=2; end
			9513: begin bcd3<=9;bcd2<=5;bcd1<=1;bcd0<=3; end
			9514: begin bcd3<=9;bcd2<=5;bcd1<=1;bcd0<=4; end
			9515: begin bcd3<=9;bcd2<=5;bcd1<=1;bcd0<=5; end
			9516: begin bcd3<=9;bcd2<=5;bcd1<=1;bcd0<=6; end
			9517: begin bcd3<=9;bcd2<=5;bcd1<=1;bcd0<=7; end
			9518: begin bcd3<=9;bcd2<=5;bcd1<=1;bcd0<=8; end
			9519: begin bcd3<=9;bcd2<=5;bcd1<=1;bcd0<=9; end
			9520: begin bcd3<=9;bcd2<=5;bcd1<=2;bcd0<=0; end
			9521: begin bcd3<=9;bcd2<=5;bcd1<=2;bcd0<=1; end
			9522: begin bcd3<=9;bcd2<=5;bcd1<=2;bcd0<=2; end
			9523: begin bcd3<=9;bcd2<=5;bcd1<=2;bcd0<=3; end
			9524: begin bcd3<=9;bcd2<=5;bcd1<=2;bcd0<=4; end
			9525: begin bcd3<=9;bcd2<=5;bcd1<=2;bcd0<=5; end
			9526: begin bcd3<=9;bcd2<=5;bcd1<=2;bcd0<=6; end
			9527: begin bcd3<=9;bcd2<=5;bcd1<=2;bcd0<=7; end
			9528: begin bcd3<=9;bcd2<=5;bcd1<=2;bcd0<=8; end
			9529: begin bcd3<=9;bcd2<=5;bcd1<=2;bcd0<=9; end
			9530: begin bcd3<=9;bcd2<=5;bcd1<=3;bcd0<=0; end
			9531: begin bcd3<=9;bcd2<=5;bcd1<=3;bcd0<=1; end
			9532: begin bcd3<=9;bcd2<=5;bcd1<=3;bcd0<=2; end
			9533: begin bcd3<=9;bcd2<=5;bcd1<=3;bcd0<=3; end
			9534: begin bcd3<=9;bcd2<=5;bcd1<=3;bcd0<=4; end
			9535: begin bcd3<=9;bcd2<=5;bcd1<=3;bcd0<=5; end
			9536: begin bcd3<=9;bcd2<=5;bcd1<=3;bcd0<=6; end
			9537: begin bcd3<=9;bcd2<=5;bcd1<=3;bcd0<=7; end
			9538: begin bcd3<=9;bcd2<=5;bcd1<=3;bcd0<=8; end
			9539: begin bcd3<=9;bcd2<=5;bcd1<=3;bcd0<=9; end
			9540: begin bcd3<=9;bcd2<=5;bcd1<=4;bcd0<=0; end
			9541: begin bcd3<=9;bcd2<=5;bcd1<=4;bcd0<=1; end
			9542: begin bcd3<=9;bcd2<=5;bcd1<=4;bcd0<=2; end
			9543: begin bcd3<=9;bcd2<=5;bcd1<=4;bcd0<=3; end
			9544: begin bcd3<=9;bcd2<=5;bcd1<=4;bcd0<=4; end
			9545: begin bcd3<=9;bcd2<=5;bcd1<=4;bcd0<=5; end
			9546: begin bcd3<=9;bcd2<=5;bcd1<=4;bcd0<=6; end
			9547: begin bcd3<=9;bcd2<=5;bcd1<=4;bcd0<=7; end
			9548: begin bcd3<=9;bcd2<=5;bcd1<=4;bcd0<=8; end
			9549: begin bcd3<=9;bcd2<=5;bcd1<=4;bcd0<=9; end
			9550: begin bcd3<=9;bcd2<=5;bcd1<=5;bcd0<=0; end
			9551: begin bcd3<=9;bcd2<=5;bcd1<=5;bcd0<=1; end
			9552: begin bcd3<=9;bcd2<=5;bcd1<=5;bcd0<=2; end
			9553: begin bcd3<=9;bcd2<=5;bcd1<=5;bcd0<=3; end
			9554: begin bcd3<=9;bcd2<=5;bcd1<=5;bcd0<=4; end
			9555: begin bcd3<=9;bcd2<=5;bcd1<=5;bcd0<=5; end
			9556: begin bcd3<=9;bcd2<=5;bcd1<=5;bcd0<=6; end
			9557: begin bcd3<=9;bcd2<=5;bcd1<=5;bcd0<=7; end
			9558: begin bcd3<=9;bcd2<=5;bcd1<=5;bcd0<=8; end
			9559: begin bcd3<=9;bcd2<=5;bcd1<=5;bcd0<=9; end
			9560: begin bcd3<=9;bcd2<=5;bcd1<=6;bcd0<=0; end
			9561: begin bcd3<=9;bcd2<=5;bcd1<=6;bcd0<=1; end
			9562: begin bcd3<=9;bcd2<=5;bcd1<=6;bcd0<=2; end
			9563: begin bcd3<=9;bcd2<=5;bcd1<=6;bcd0<=3; end
			9564: begin bcd3<=9;bcd2<=5;bcd1<=6;bcd0<=4; end
			9565: begin bcd3<=9;bcd2<=5;bcd1<=6;bcd0<=5; end
			9566: begin bcd3<=9;bcd2<=5;bcd1<=6;bcd0<=6; end
			9567: begin bcd3<=9;bcd2<=5;bcd1<=6;bcd0<=7; end
			9568: begin bcd3<=9;bcd2<=5;bcd1<=6;bcd0<=8; end
			9569: begin bcd3<=9;bcd2<=5;bcd1<=6;bcd0<=9; end
			9570: begin bcd3<=9;bcd2<=5;bcd1<=7;bcd0<=0; end
			9571: begin bcd3<=9;bcd2<=5;bcd1<=7;bcd0<=1; end
			9572: begin bcd3<=9;bcd2<=5;bcd1<=7;bcd0<=2; end
			9573: begin bcd3<=9;bcd2<=5;bcd1<=7;bcd0<=3; end
			9574: begin bcd3<=9;bcd2<=5;bcd1<=7;bcd0<=4; end
			9575: begin bcd3<=9;bcd2<=5;bcd1<=7;bcd0<=5; end
			9576: begin bcd3<=9;bcd2<=5;bcd1<=7;bcd0<=6; end
			9577: begin bcd3<=9;bcd2<=5;bcd1<=7;bcd0<=7; end
			9578: begin bcd3<=9;bcd2<=5;bcd1<=7;bcd0<=8; end
			9579: begin bcd3<=9;bcd2<=5;bcd1<=7;bcd0<=9; end
			9580: begin bcd3<=9;bcd2<=5;bcd1<=8;bcd0<=0; end
			9581: begin bcd3<=9;bcd2<=5;bcd1<=8;bcd0<=1; end
			9582: begin bcd3<=9;bcd2<=5;bcd1<=8;bcd0<=2; end
			9583: begin bcd3<=9;bcd2<=5;bcd1<=8;bcd0<=3; end
			9584: begin bcd3<=9;bcd2<=5;bcd1<=8;bcd0<=4; end
			9585: begin bcd3<=9;bcd2<=5;bcd1<=8;bcd0<=5; end
			9586: begin bcd3<=9;bcd2<=5;bcd1<=8;bcd0<=6; end
			9587: begin bcd3<=9;bcd2<=5;bcd1<=8;bcd0<=7; end
			9588: begin bcd3<=9;bcd2<=5;bcd1<=8;bcd0<=8; end
			9589: begin bcd3<=9;bcd2<=5;bcd1<=8;bcd0<=9; end
			9590: begin bcd3<=9;bcd2<=5;bcd1<=9;bcd0<=0; end
			9591: begin bcd3<=9;bcd2<=5;bcd1<=9;bcd0<=1; end
			9592: begin bcd3<=9;bcd2<=5;bcd1<=9;bcd0<=2; end
			9593: begin bcd3<=9;bcd2<=5;bcd1<=9;bcd0<=3; end
			9594: begin bcd3<=9;bcd2<=5;bcd1<=9;bcd0<=4; end
			9595: begin bcd3<=9;bcd2<=5;bcd1<=9;bcd0<=5; end
			9596: begin bcd3<=9;bcd2<=5;bcd1<=9;bcd0<=6; end
			9597: begin bcd3<=9;bcd2<=5;bcd1<=9;bcd0<=7; end
			9598: begin bcd3<=9;bcd2<=5;bcd1<=9;bcd0<=8; end
			9599: begin bcd3<=9;bcd2<=5;bcd1<=9;bcd0<=9; end
			9600: begin bcd3<=9;bcd2<=6;bcd1<=0;bcd0<=0; end
			9601: begin bcd3<=9;bcd2<=6;bcd1<=0;bcd0<=1; end
			9602: begin bcd3<=9;bcd2<=6;bcd1<=0;bcd0<=2; end
			9603: begin bcd3<=9;bcd2<=6;bcd1<=0;bcd0<=3; end
			9604: begin bcd3<=9;bcd2<=6;bcd1<=0;bcd0<=4; end
			9605: begin bcd3<=9;bcd2<=6;bcd1<=0;bcd0<=5; end
			9606: begin bcd3<=9;bcd2<=6;bcd1<=0;bcd0<=6; end
			9607: begin bcd3<=9;bcd2<=6;bcd1<=0;bcd0<=7; end
			9608: begin bcd3<=9;bcd2<=6;bcd1<=0;bcd0<=8; end
			9609: begin bcd3<=9;bcd2<=6;bcd1<=0;bcd0<=9; end
			9610: begin bcd3<=9;bcd2<=6;bcd1<=1;bcd0<=0; end
			9611: begin bcd3<=9;bcd2<=6;bcd1<=1;bcd0<=1; end
			9612: begin bcd3<=9;bcd2<=6;bcd1<=1;bcd0<=2; end
			9613: begin bcd3<=9;bcd2<=6;bcd1<=1;bcd0<=3; end
			9614: begin bcd3<=9;bcd2<=6;bcd1<=1;bcd0<=4; end
			9615: begin bcd3<=9;bcd2<=6;bcd1<=1;bcd0<=5; end
			9616: begin bcd3<=9;bcd2<=6;bcd1<=1;bcd0<=6; end
			9617: begin bcd3<=9;bcd2<=6;bcd1<=1;bcd0<=7; end
			9618: begin bcd3<=9;bcd2<=6;bcd1<=1;bcd0<=8; end
			9619: begin bcd3<=9;bcd2<=6;bcd1<=1;bcd0<=9; end
			9620: begin bcd3<=9;bcd2<=6;bcd1<=2;bcd0<=0; end
			9621: begin bcd3<=9;bcd2<=6;bcd1<=2;bcd0<=1; end
			9622: begin bcd3<=9;bcd2<=6;bcd1<=2;bcd0<=2; end
			9623: begin bcd3<=9;bcd2<=6;bcd1<=2;bcd0<=3; end
			9624: begin bcd3<=9;bcd2<=6;bcd1<=2;bcd0<=4; end
			9625: begin bcd3<=9;bcd2<=6;bcd1<=2;bcd0<=5; end
			9626: begin bcd3<=9;bcd2<=6;bcd1<=2;bcd0<=6; end
			9627: begin bcd3<=9;bcd2<=6;bcd1<=2;bcd0<=7; end
			9628: begin bcd3<=9;bcd2<=6;bcd1<=2;bcd0<=8; end
			9629: begin bcd3<=9;bcd2<=6;bcd1<=2;bcd0<=9; end
			9630: begin bcd3<=9;bcd2<=6;bcd1<=3;bcd0<=0; end
			9631: begin bcd3<=9;bcd2<=6;bcd1<=3;bcd0<=1; end
			9632: begin bcd3<=9;bcd2<=6;bcd1<=3;bcd0<=2; end
			9633: begin bcd3<=9;bcd2<=6;bcd1<=3;bcd0<=3; end
			9634: begin bcd3<=9;bcd2<=6;bcd1<=3;bcd0<=4; end
			9635: begin bcd3<=9;bcd2<=6;bcd1<=3;bcd0<=5; end
			9636: begin bcd3<=9;bcd2<=6;bcd1<=3;bcd0<=6; end
			9637: begin bcd3<=9;bcd2<=6;bcd1<=3;bcd0<=7; end
			9638: begin bcd3<=9;bcd2<=6;bcd1<=3;bcd0<=8; end
			9639: begin bcd3<=9;bcd2<=6;bcd1<=3;bcd0<=9; end
			9640: begin bcd3<=9;bcd2<=6;bcd1<=4;bcd0<=0; end
			9641: begin bcd3<=9;bcd2<=6;bcd1<=4;bcd0<=1; end
			9642: begin bcd3<=9;bcd2<=6;bcd1<=4;bcd0<=2; end
			9643: begin bcd3<=9;bcd2<=6;bcd1<=4;bcd0<=3; end
			9644: begin bcd3<=9;bcd2<=6;bcd1<=4;bcd0<=4; end
			9645: begin bcd3<=9;bcd2<=6;bcd1<=4;bcd0<=5; end
			9646: begin bcd3<=9;bcd2<=6;bcd1<=4;bcd0<=6; end
			9647: begin bcd3<=9;bcd2<=6;bcd1<=4;bcd0<=7; end
			9648: begin bcd3<=9;bcd2<=6;bcd1<=4;bcd0<=8; end
			9649: begin bcd3<=9;bcd2<=6;bcd1<=4;bcd0<=9; end
			9650: begin bcd3<=9;bcd2<=6;bcd1<=5;bcd0<=0; end
			9651: begin bcd3<=9;bcd2<=6;bcd1<=5;bcd0<=1; end
			9652: begin bcd3<=9;bcd2<=6;bcd1<=5;bcd0<=2; end
			9653: begin bcd3<=9;bcd2<=6;bcd1<=5;bcd0<=3; end
			9654: begin bcd3<=9;bcd2<=6;bcd1<=5;bcd0<=4; end
			9655: begin bcd3<=9;bcd2<=6;bcd1<=5;bcd0<=5; end
			9656: begin bcd3<=9;bcd2<=6;bcd1<=5;bcd0<=6; end
			9657: begin bcd3<=9;bcd2<=6;bcd1<=5;bcd0<=7; end
			9658: begin bcd3<=9;bcd2<=6;bcd1<=5;bcd0<=8; end
			9659: begin bcd3<=9;bcd2<=6;bcd1<=5;bcd0<=9; end
			9660: begin bcd3<=9;bcd2<=6;bcd1<=6;bcd0<=0; end
			9661: begin bcd3<=9;bcd2<=6;bcd1<=6;bcd0<=1; end
			9662: begin bcd3<=9;bcd2<=6;bcd1<=6;bcd0<=2; end
			9663: begin bcd3<=9;bcd2<=6;bcd1<=6;bcd0<=3; end
			9664: begin bcd3<=9;bcd2<=6;bcd1<=6;bcd0<=4; end
			9665: begin bcd3<=9;bcd2<=6;bcd1<=6;bcd0<=5; end
			9666: begin bcd3<=9;bcd2<=6;bcd1<=6;bcd0<=6; end
			9667: begin bcd3<=9;bcd2<=6;bcd1<=6;bcd0<=7; end
			9668: begin bcd3<=9;bcd2<=6;bcd1<=6;bcd0<=8; end
			9669: begin bcd3<=9;bcd2<=6;bcd1<=6;bcd0<=9; end
			9670: begin bcd3<=9;bcd2<=6;bcd1<=7;bcd0<=0; end
			9671: begin bcd3<=9;bcd2<=6;bcd1<=7;bcd0<=1; end
			9672: begin bcd3<=9;bcd2<=6;bcd1<=7;bcd0<=2; end
			9673: begin bcd3<=9;bcd2<=6;bcd1<=7;bcd0<=3; end
			9674: begin bcd3<=9;bcd2<=6;bcd1<=7;bcd0<=4; end
			9675: begin bcd3<=9;bcd2<=6;bcd1<=7;bcd0<=5; end
			9676: begin bcd3<=9;bcd2<=6;bcd1<=7;bcd0<=6; end
			9677: begin bcd3<=9;bcd2<=6;bcd1<=7;bcd0<=7; end
			9678: begin bcd3<=9;bcd2<=6;bcd1<=7;bcd0<=8; end
			9679: begin bcd3<=9;bcd2<=6;bcd1<=7;bcd0<=9; end
			9680: begin bcd3<=9;bcd2<=6;bcd1<=8;bcd0<=0; end
			9681: begin bcd3<=9;bcd2<=6;bcd1<=8;bcd0<=1; end
			9682: begin bcd3<=9;bcd2<=6;bcd1<=8;bcd0<=2; end
			9683: begin bcd3<=9;bcd2<=6;bcd1<=8;bcd0<=3; end
			9684: begin bcd3<=9;bcd2<=6;bcd1<=8;bcd0<=4; end
			9685: begin bcd3<=9;bcd2<=6;bcd1<=8;bcd0<=5; end
			9686: begin bcd3<=9;bcd2<=6;bcd1<=8;bcd0<=6; end
			9687: begin bcd3<=9;bcd2<=6;bcd1<=8;bcd0<=7; end
			9688: begin bcd3<=9;bcd2<=6;bcd1<=8;bcd0<=8; end
			9689: begin bcd3<=9;bcd2<=6;bcd1<=8;bcd0<=9; end
			9690: begin bcd3<=9;bcd2<=6;bcd1<=9;bcd0<=0; end
			9691: begin bcd3<=9;bcd2<=6;bcd1<=9;bcd0<=1; end
			9692: begin bcd3<=9;bcd2<=6;bcd1<=9;bcd0<=2; end
			9693: begin bcd3<=9;bcd2<=6;bcd1<=9;bcd0<=3; end
			9694: begin bcd3<=9;bcd2<=6;bcd1<=9;bcd0<=4; end
			9695: begin bcd3<=9;bcd2<=6;bcd1<=9;bcd0<=5; end
			9696: begin bcd3<=9;bcd2<=6;bcd1<=9;bcd0<=6; end
			9697: begin bcd3<=9;bcd2<=6;bcd1<=9;bcd0<=7; end
			9698: begin bcd3<=9;bcd2<=6;bcd1<=9;bcd0<=8; end
			9699: begin bcd3<=9;bcd2<=6;bcd1<=9;bcd0<=9; end
			9700: begin bcd3<=9;bcd2<=7;bcd1<=0;bcd0<=0; end
			9701: begin bcd3<=9;bcd2<=7;bcd1<=0;bcd0<=1; end
			9702: begin bcd3<=9;bcd2<=7;bcd1<=0;bcd0<=2; end
			9703: begin bcd3<=9;bcd2<=7;bcd1<=0;bcd0<=3; end
			9704: begin bcd3<=9;bcd2<=7;bcd1<=0;bcd0<=4; end
			9705: begin bcd3<=9;bcd2<=7;bcd1<=0;bcd0<=5; end
			9706: begin bcd3<=9;bcd2<=7;bcd1<=0;bcd0<=6; end
			9707: begin bcd3<=9;bcd2<=7;bcd1<=0;bcd0<=7; end
			9708: begin bcd3<=9;bcd2<=7;bcd1<=0;bcd0<=8; end
			9709: begin bcd3<=9;bcd2<=7;bcd1<=0;bcd0<=9; end
			9710: begin bcd3<=9;bcd2<=7;bcd1<=1;bcd0<=0; end
			9711: begin bcd3<=9;bcd2<=7;bcd1<=1;bcd0<=1; end
			9712: begin bcd3<=9;bcd2<=7;bcd1<=1;bcd0<=2; end
			9713: begin bcd3<=9;bcd2<=7;bcd1<=1;bcd0<=3; end
			9714: begin bcd3<=9;bcd2<=7;bcd1<=1;bcd0<=4; end
			9715: begin bcd3<=9;bcd2<=7;bcd1<=1;bcd0<=5; end
			9716: begin bcd3<=9;bcd2<=7;bcd1<=1;bcd0<=6; end
			9717: begin bcd3<=9;bcd2<=7;bcd1<=1;bcd0<=7; end
			9718: begin bcd3<=9;bcd2<=7;bcd1<=1;bcd0<=8; end
			9719: begin bcd3<=9;bcd2<=7;bcd1<=1;bcd0<=9; end
			9720: begin bcd3<=9;bcd2<=7;bcd1<=2;bcd0<=0; end
			9721: begin bcd3<=9;bcd2<=7;bcd1<=2;bcd0<=1; end
			9722: begin bcd3<=9;bcd2<=7;bcd1<=2;bcd0<=2; end
			9723: begin bcd3<=9;bcd2<=7;bcd1<=2;bcd0<=3; end
			9724: begin bcd3<=9;bcd2<=7;bcd1<=2;bcd0<=4; end
			9725: begin bcd3<=9;bcd2<=7;bcd1<=2;bcd0<=5; end
			9726: begin bcd3<=9;bcd2<=7;bcd1<=2;bcd0<=6; end
			9727: begin bcd3<=9;bcd2<=7;bcd1<=2;bcd0<=7; end
			9728: begin bcd3<=9;bcd2<=7;bcd1<=2;bcd0<=8; end
			9729: begin bcd3<=9;bcd2<=7;bcd1<=2;bcd0<=9; end
			9730: begin bcd3<=9;bcd2<=7;bcd1<=3;bcd0<=0; end
			9731: begin bcd3<=9;bcd2<=7;bcd1<=3;bcd0<=1; end
			9732: begin bcd3<=9;bcd2<=7;bcd1<=3;bcd0<=2; end
			9733: begin bcd3<=9;bcd2<=7;bcd1<=3;bcd0<=3; end
			9734: begin bcd3<=9;bcd2<=7;bcd1<=3;bcd0<=4; end
			9735: begin bcd3<=9;bcd2<=7;bcd1<=3;bcd0<=5; end
			9736: begin bcd3<=9;bcd2<=7;bcd1<=3;bcd0<=6; end
			9737: begin bcd3<=9;bcd2<=7;bcd1<=3;bcd0<=7; end
			9738: begin bcd3<=9;bcd2<=7;bcd1<=3;bcd0<=8; end
			9739: begin bcd3<=9;bcd2<=7;bcd1<=3;bcd0<=9; end
			9740: begin bcd3<=9;bcd2<=7;bcd1<=4;bcd0<=0; end
			9741: begin bcd3<=9;bcd2<=7;bcd1<=4;bcd0<=1; end
			9742: begin bcd3<=9;bcd2<=7;bcd1<=4;bcd0<=2; end
			9743: begin bcd3<=9;bcd2<=7;bcd1<=4;bcd0<=3; end
			9744: begin bcd3<=9;bcd2<=7;bcd1<=4;bcd0<=4; end
			9745: begin bcd3<=9;bcd2<=7;bcd1<=4;bcd0<=5; end
			9746: begin bcd3<=9;bcd2<=7;bcd1<=4;bcd0<=6; end
			9747: begin bcd3<=9;bcd2<=7;bcd1<=4;bcd0<=7; end
			9748: begin bcd3<=9;bcd2<=7;bcd1<=4;bcd0<=8; end
			9749: begin bcd3<=9;bcd2<=7;bcd1<=4;bcd0<=9; end
			9750: begin bcd3<=9;bcd2<=7;bcd1<=5;bcd0<=0; end
			9751: begin bcd3<=9;bcd2<=7;bcd1<=5;bcd0<=1; end
			9752: begin bcd3<=9;bcd2<=7;bcd1<=5;bcd0<=2; end
			9753: begin bcd3<=9;bcd2<=7;bcd1<=5;bcd0<=3; end
			9754: begin bcd3<=9;bcd2<=7;bcd1<=5;bcd0<=4; end
			9755: begin bcd3<=9;bcd2<=7;bcd1<=5;bcd0<=5; end
			9756: begin bcd3<=9;bcd2<=7;bcd1<=5;bcd0<=6; end
			9757: begin bcd3<=9;bcd2<=7;bcd1<=5;bcd0<=7; end
			9758: begin bcd3<=9;bcd2<=7;bcd1<=5;bcd0<=8; end
			9759: begin bcd3<=9;bcd2<=7;bcd1<=5;bcd0<=9; end
			9760: begin bcd3<=9;bcd2<=7;bcd1<=6;bcd0<=0; end
			9761: begin bcd3<=9;bcd2<=7;bcd1<=6;bcd0<=1; end
			9762: begin bcd3<=9;bcd2<=7;bcd1<=6;bcd0<=2; end
			9763: begin bcd3<=9;bcd2<=7;bcd1<=6;bcd0<=3; end
			9764: begin bcd3<=9;bcd2<=7;bcd1<=6;bcd0<=4; end
			9765: begin bcd3<=9;bcd2<=7;bcd1<=6;bcd0<=5; end
			9766: begin bcd3<=9;bcd2<=7;bcd1<=6;bcd0<=6; end
			9767: begin bcd3<=9;bcd2<=7;bcd1<=6;bcd0<=7; end
			9768: begin bcd3<=9;bcd2<=7;bcd1<=6;bcd0<=8; end
			9769: begin bcd3<=9;bcd2<=7;bcd1<=6;bcd0<=9; end
			9770: begin bcd3<=9;bcd2<=7;bcd1<=7;bcd0<=0; end
			9771: begin bcd3<=9;bcd2<=7;bcd1<=7;bcd0<=1; end
			9772: begin bcd3<=9;bcd2<=7;bcd1<=7;bcd0<=2; end
			9773: begin bcd3<=9;bcd2<=7;bcd1<=7;bcd0<=3; end
			9774: begin bcd3<=9;bcd2<=7;bcd1<=7;bcd0<=4; end
			9775: begin bcd3<=9;bcd2<=7;bcd1<=7;bcd0<=5; end
			9776: begin bcd3<=9;bcd2<=7;bcd1<=7;bcd0<=6; end
			9777: begin bcd3<=9;bcd2<=7;bcd1<=7;bcd0<=7; end
			9778: begin bcd3<=9;bcd2<=7;bcd1<=7;bcd0<=8; end
			9779: begin bcd3<=9;bcd2<=7;bcd1<=7;bcd0<=9; end
			9780: begin bcd3<=9;bcd2<=7;bcd1<=8;bcd0<=0; end
			9781: begin bcd3<=9;bcd2<=7;bcd1<=8;bcd0<=1; end
			9782: begin bcd3<=9;bcd2<=7;bcd1<=8;bcd0<=2; end
			9783: begin bcd3<=9;bcd2<=7;bcd1<=8;bcd0<=3; end
			9784: begin bcd3<=9;bcd2<=7;bcd1<=8;bcd0<=4; end
			9785: begin bcd3<=9;bcd2<=7;bcd1<=8;bcd0<=5; end
			9786: begin bcd3<=9;bcd2<=7;bcd1<=8;bcd0<=6; end
			9787: begin bcd3<=9;bcd2<=7;bcd1<=8;bcd0<=7; end
			9788: begin bcd3<=9;bcd2<=7;bcd1<=8;bcd0<=8; end
			9789: begin bcd3<=9;bcd2<=7;bcd1<=8;bcd0<=9; end
			9790: begin bcd3<=9;bcd2<=7;bcd1<=9;bcd0<=0; end
			9791: begin bcd3<=9;bcd2<=7;bcd1<=9;bcd0<=1; end
			9792: begin bcd3<=9;bcd2<=7;bcd1<=9;bcd0<=2; end
			9793: begin bcd3<=9;bcd2<=7;bcd1<=9;bcd0<=3; end
			9794: begin bcd3<=9;bcd2<=7;bcd1<=9;bcd0<=4; end
			9795: begin bcd3<=9;bcd2<=7;bcd1<=9;bcd0<=5; end
			9796: begin bcd3<=9;bcd2<=7;bcd1<=9;bcd0<=6; end
			9797: begin bcd3<=9;bcd2<=7;bcd1<=9;bcd0<=7; end
			9798: begin bcd3<=9;bcd2<=7;bcd1<=9;bcd0<=8; end
			9799: begin bcd3<=9;bcd2<=7;bcd1<=9;bcd0<=9; end
			9800: begin bcd3<=9;bcd2<=8;bcd1<=0;bcd0<=0; end
			9801: begin bcd3<=9;bcd2<=8;bcd1<=0;bcd0<=1; end
			9802: begin bcd3<=9;bcd2<=8;bcd1<=0;bcd0<=2; end
			9803: begin bcd3<=9;bcd2<=8;bcd1<=0;bcd0<=3; end
			9804: begin bcd3<=9;bcd2<=8;bcd1<=0;bcd0<=4; end
			9805: begin bcd3<=9;bcd2<=8;bcd1<=0;bcd0<=5; end
			9806: begin bcd3<=9;bcd2<=8;bcd1<=0;bcd0<=6; end
			9807: begin bcd3<=9;bcd2<=8;bcd1<=0;bcd0<=7; end
			9808: begin bcd3<=9;bcd2<=8;bcd1<=0;bcd0<=8; end
			9809: begin bcd3<=9;bcd2<=8;bcd1<=0;bcd0<=9; end
			9810: begin bcd3<=9;bcd2<=8;bcd1<=1;bcd0<=0; end
			9811: begin bcd3<=9;bcd2<=8;bcd1<=1;bcd0<=1; end
			9812: begin bcd3<=9;bcd2<=8;bcd1<=1;bcd0<=2; end
			9813: begin bcd3<=9;bcd2<=8;bcd1<=1;bcd0<=3; end
			9814: begin bcd3<=9;bcd2<=8;bcd1<=1;bcd0<=4; end
			9815: begin bcd3<=9;bcd2<=8;bcd1<=1;bcd0<=5; end
			9816: begin bcd3<=9;bcd2<=8;bcd1<=1;bcd0<=6; end
			9817: begin bcd3<=9;bcd2<=8;bcd1<=1;bcd0<=7; end
			9818: begin bcd3<=9;bcd2<=8;bcd1<=1;bcd0<=8; end
			9819: begin bcd3<=9;bcd2<=8;bcd1<=1;bcd0<=9; end
			9820: begin bcd3<=9;bcd2<=8;bcd1<=2;bcd0<=0; end
			9821: begin bcd3<=9;bcd2<=8;bcd1<=2;bcd0<=1; end
			9822: begin bcd3<=9;bcd2<=8;bcd1<=2;bcd0<=2; end
			9823: begin bcd3<=9;bcd2<=8;bcd1<=2;bcd0<=3; end
			9824: begin bcd3<=9;bcd2<=8;bcd1<=2;bcd0<=4; end
			9825: begin bcd3<=9;bcd2<=8;bcd1<=2;bcd0<=5; end
			9826: begin bcd3<=9;bcd2<=8;bcd1<=2;bcd0<=6; end
			9827: begin bcd3<=9;bcd2<=8;bcd1<=2;bcd0<=7; end
			9828: begin bcd3<=9;bcd2<=8;bcd1<=2;bcd0<=8; end
			9829: begin bcd3<=9;bcd2<=8;bcd1<=2;bcd0<=9; end
			9830: begin bcd3<=9;bcd2<=8;bcd1<=3;bcd0<=0; end
			9831: begin bcd3<=9;bcd2<=8;bcd1<=3;bcd0<=1; end
			9832: begin bcd3<=9;bcd2<=8;bcd1<=3;bcd0<=2; end
			9833: begin bcd3<=9;bcd2<=8;bcd1<=3;bcd0<=3; end
			9834: begin bcd3<=9;bcd2<=8;bcd1<=3;bcd0<=4; end
			9835: begin bcd3<=9;bcd2<=8;bcd1<=3;bcd0<=5; end
			9836: begin bcd3<=9;bcd2<=8;bcd1<=3;bcd0<=6; end
			9837: begin bcd3<=9;bcd2<=8;bcd1<=3;bcd0<=7; end
			9838: begin bcd3<=9;bcd2<=8;bcd1<=3;bcd0<=8; end
			9839: begin bcd3<=9;bcd2<=8;bcd1<=3;bcd0<=9; end
			9840: begin bcd3<=9;bcd2<=8;bcd1<=4;bcd0<=0; end
			9841: begin bcd3<=9;bcd2<=8;bcd1<=4;bcd0<=1; end
			9842: begin bcd3<=9;bcd2<=8;bcd1<=4;bcd0<=2; end
			9843: begin bcd3<=9;bcd2<=8;bcd1<=4;bcd0<=3; end
			9844: begin bcd3<=9;bcd2<=8;bcd1<=4;bcd0<=4; end
			9845: begin bcd3<=9;bcd2<=8;bcd1<=4;bcd0<=5; end
			9846: begin bcd3<=9;bcd2<=8;bcd1<=4;bcd0<=6; end
			9847: begin bcd3<=9;bcd2<=8;bcd1<=4;bcd0<=7; end
			9848: begin bcd3<=9;bcd2<=8;bcd1<=4;bcd0<=8; end
			9849: begin bcd3<=9;bcd2<=8;bcd1<=4;bcd0<=9; end
			9850: begin bcd3<=9;bcd2<=8;bcd1<=5;bcd0<=0; end
			9851: begin bcd3<=9;bcd2<=8;bcd1<=5;bcd0<=1; end
			9852: begin bcd3<=9;bcd2<=8;bcd1<=5;bcd0<=2; end
			9853: begin bcd3<=9;bcd2<=8;bcd1<=5;bcd0<=3; end
			9854: begin bcd3<=9;bcd2<=8;bcd1<=5;bcd0<=4; end
			9855: begin bcd3<=9;bcd2<=8;bcd1<=5;bcd0<=5; end
			9856: begin bcd3<=9;bcd2<=8;bcd1<=5;bcd0<=6; end
			9857: begin bcd3<=9;bcd2<=8;bcd1<=5;bcd0<=7; end
			9858: begin bcd3<=9;bcd2<=8;bcd1<=5;bcd0<=8; end
			9859: begin bcd3<=9;bcd2<=8;bcd1<=5;bcd0<=9; end
			9860: begin bcd3<=9;bcd2<=8;bcd1<=6;bcd0<=0; end
			9861: begin bcd3<=9;bcd2<=8;bcd1<=6;bcd0<=1; end
			9862: begin bcd3<=9;bcd2<=8;bcd1<=6;bcd0<=2; end
			9863: begin bcd3<=9;bcd2<=8;bcd1<=6;bcd0<=3; end
			9864: begin bcd3<=9;bcd2<=8;bcd1<=6;bcd0<=4; end
			9865: begin bcd3<=9;bcd2<=8;bcd1<=6;bcd0<=5; end
			9866: begin bcd3<=9;bcd2<=8;bcd1<=6;bcd0<=6; end
			9867: begin bcd3<=9;bcd2<=8;bcd1<=6;bcd0<=7; end
			9868: begin bcd3<=9;bcd2<=8;bcd1<=6;bcd0<=8; end
			9869: begin bcd3<=9;bcd2<=8;bcd1<=6;bcd0<=9; end
			9870: begin bcd3<=9;bcd2<=8;bcd1<=7;bcd0<=0; end
			9871: begin bcd3<=9;bcd2<=8;bcd1<=7;bcd0<=1; end
			9872: begin bcd3<=9;bcd2<=8;bcd1<=7;bcd0<=2; end
			9873: begin bcd3<=9;bcd2<=8;bcd1<=7;bcd0<=3; end
			9874: begin bcd3<=9;bcd2<=8;bcd1<=7;bcd0<=4; end
			9875: begin bcd3<=9;bcd2<=8;bcd1<=7;bcd0<=5; end
			9876: begin bcd3<=9;bcd2<=8;bcd1<=7;bcd0<=6; end
			9877: begin bcd3<=9;bcd2<=8;bcd1<=7;bcd0<=7; end
			9878: begin bcd3<=9;bcd2<=8;bcd1<=7;bcd0<=8; end
			9879: begin bcd3<=9;bcd2<=8;bcd1<=7;bcd0<=9; end
			9880: begin bcd3<=9;bcd2<=8;bcd1<=8;bcd0<=0; end
			9881: begin bcd3<=9;bcd2<=8;bcd1<=8;bcd0<=1; end
			9882: begin bcd3<=9;bcd2<=8;bcd1<=8;bcd0<=2; end
			9883: begin bcd3<=9;bcd2<=8;bcd1<=8;bcd0<=3; end
			9884: begin bcd3<=9;bcd2<=8;bcd1<=8;bcd0<=4; end
			9885: begin bcd3<=9;bcd2<=8;bcd1<=8;bcd0<=5; end
			9886: begin bcd3<=9;bcd2<=8;bcd1<=8;bcd0<=6; end
			9887: begin bcd3<=9;bcd2<=8;bcd1<=8;bcd0<=7; end
			9888: begin bcd3<=9;bcd2<=8;bcd1<=8;bcd0<=8; end
			9889: begin bcd3<=9;bcd2<=8;bcd1<=8;bcd0<=9; end
			9890: begin bcd3<=9;bcd2<=8;bcd1<=9;bcd0<=0; end
			9891: begin bcd3<=9;bcd2<=8;bcd1<=9;bcd0<=1; end
			9892: begin bcd3<=9;bcd2<=8;bcd1<=9;bcd0<=2; end
			9893: begin bcd3<=9;bcd2<=8;bcd1<=9;bcd0<=3; end
			9894: begin bcd3<=9;bcd2<=8;bcd1<=9;bcd0<=4; end
			9895: begin bcd3<=9;bcd2<=8;bcd1<=9;bcd0<=5; end
			9896: begin bcd3<=9;bcd2<=8;bcd1<=9;bcd0<=6; end
			9897: begin bcd3<=9;bcd2<=8;bcd1<=9;bcd0<=7; end
			9898: begin bcd3<=9;bcd2<=8;bcd1<=9;bcd0<=8; end
			9899: begin bcd3<=9;bcd2<=8;bcd1<=9;bcd0<=9; end
			9900: begin bcd3<=9;bcd2<=9;bcd1<=0;bcd0<=0; end
			9901: begin bcd3<=9;bcd2<=9;bcd1<=0;bcd0<=1; end
			9902: begin bcd3<=9;bcd2<=9;bcd1<=0;bcd0<=2; end
			9903: begin bcd3<=9;bcd2<=9;bcd1<=0;bcd0<=3; end
			9904: begin bcd3<=9;bcd2<=9;bcd1<=0;bcd0<=4; end
			9905: begin bcd3<=9;bcd2<=9;bcd1<=0;bcd0<=5; end
			9906: begin bcd3<=9;bcd2<=9;bcd1<=0;bcd0<=6; end
			9907: begin bcd3<=9;bcd2<=9;bcd1<=0;bcd0<=7; end
			9908: begin bcd3<=9;bcd2<=9;bcd1<=0;bcd0<=8; end
			9909: begin bcd3<=9;bcd2<=9;bcd1<=0;bcd0<=9; end
			9910: begin bcd3<=9;bcd2<=9;bcd1<=1;bcd0<=0; end
			9911: begin bcd3<=9;bcd2<=9;bcd1<=1;bcd0<=1; end
			9912: begin bcd3<=9;bcd2<=9;bcd1<=1;bcd0<=2; end
			9913: begin bcd3<=9;bcd2<=9;bcd1<=1;bcd0<=3; end
			9914: begin bcd3<=9;bcd2<=9;bcd1<=1;bcd0<=4; end
			9915: begin bcd3<=9;bcd2<=9;bcd1<=1;bcd0<=5; end
			9916: begin bcd3<=9;bcd2<=9;bcd1<=1;bcd0<=6; end
			9917: begin bcd3<=9;bcd2<=9;bcd1<=1;bcd0<=7; end
			9918: begin bcd3<=9;bcd2<=9;bcd1<=1;bcd0<=8; end
			9919: begin bcd3<=9;bcd2<=9;bcd1<=1;bcd0<=9; end
			9920: begin bcd3<=9;bcd2<=9;bcd1<=2;bcd0<=0; end
			9921: begin bcd3<=9;bcd2<=9;bcd1<=2;bcd0<=1; end
			9922: begin bcd3<=9;bcd2<=9;bcd1<=2;bcd0<=2; end
			9923: begin bcd3<=9;bcd2<=9;bcd1<=2;bcd0<=3; end
			9924: begin bcd3<=9;bcd2<=9;bcd1<=2;bcd0<=4; end
			9925: begin bcd3<=9;bcd2<=9;bcd1<=2;bcd0<=5; end
			9926: begin bcd3<=9;bcd2<=9;bcd1<=2;bcd0<=6; end
			9927: begin bcd3<=9;bcd2<=9;bcd1<=2;bcd0<=7; end
			9928: begin bcd3<=9;bcd2<=9;bcd1<=2;bcd0<=8; end
			9929: begin bcd3<=9;bcd2<=9;bcd1<=2;bcd0<=9; end
			9930: begin bcd3<=9;bcd2<=9;bcd1<=3;bcd0<=0; end
			9931: begin bcd3<=9;bcd2<=9;bcd1<=3;bcd0<=1; end
			9932: begin bcd3<=9;bcd2<=9;bcd1<=3;bcd0<=2; end
			9933: begin bcd3<=9;bcd2<=9;bcd1<=3;bcd0<=3; end
			9934: begin bcd3<=9;bcd2<=9;bcd1<=3;bcd0<=4; end
			9935: begin bcd3<=9;bcd2<=9;bcd1<=3;bcd0<=5; end
			9936: begin bcd3<=9;bcd2<=9;bcd1<=3;bcd0<=6; end
			9937: begin bcd3<=9;bcd2<=9;bcd1<=3;bcd0<=7; end
			9938: begin bcd3<=9;bcd2<=9;bcd1<=3;bcd0<=8; end
			9939: begin bcd3<=9;bcd2<=9;bcd1<=3;bcd0<=9; end
			9940: begin bcd3<=9;bcd2<=9;bcd1<=4;bcd0<=0; end
			9941: begin bcd3<=9;bcd2<=9;bcd1<=4;bcd0<=1; end
			9942: begin bcd3<=9;bcd2<=9;bcd1<=4;bcd0<=2; end
			9943: begin bcd3<=9;bcd2<=9;bcd1<=4;bcd0<=3; end
			9944: begin bcd3<=9;bcd2<=9;bcd1<=4;bcd0<=4; end
			9945: begin bcd3<=9;bcd2<=9;bcd1<=4;bcd0<=5; end
			9946: begin bcd3<=9;bcd2<=9;bcd1<=4;bcd0<=6; end
			9947: begin bcd3<=9;bcd2<=9;bcd1<=4;bcd0<=7; end
			9948: begin bcd3<=9;bcd2<=9;bcd1<=4;bcd0<=8; end
			9949: begin bcd3<=9;bcd2<=9;bcd1<=4;bcd0<=9; end
			9950: begin bcd3<=9;bcd2<=9;bcd1<=5;bcd0<=0; end
			9951: begin bcd3<=9;bcd2<=9;bcd1<=5;bcd0<=1; end
			9952: begin bcd3<=9;bcd2<=9;bcd1<=5;bcd0<=2; end
			9953: begin bcd3<=9;bcd2<=9;bcd1<=5;bcd0<=3; end
			9954: begin bcd3<=9;bcd2<=9;bcd1<=5;bcd0<=4; end
			9955: begin bcd3<=9;bcd2<=9;bcd1<=5;bcd0<=5; end
			9956: begin bcd3<=9;bcd2<=9;bcd1<=5;bcd0<=6; end
			9957: begin bcd3<=9;bcd2<=9;bcd1<=5;bcd0<=7; end
			9958: begin bcd3<=9;bcd2<=9;bcd1<=5;bcd0<=8; end
			9959: begin bcd3<=9;bcd2<=9;bcd1<=5;bcd0<=9; end
			9960: begin bcd3<=9;bcd2<=9;bcd1<=6;bcd0<=0; end
			9961: begin bcd3<=9;bcd2<=9;bcd1<=6;bcd0<=1; end
			9962: begin bcd3<=9;bcd2<=9;bcd1<=6;bcd0<=2; end
			9963: begin bcd3<=9;bcd2<=9;bcd1<=6;bcd0<=3; end
			9964: begin bcd3<=9;bcd2<=9;bcd1<=6;bcd0<=4; end
			9965: begin bcd3<=9;bcd2<=9;bcd1<=6;bcd0<=5; end
			9966: begin bcd3<=9;bcd2<=9;bcd1<=6;bcd0<=6; end
			9967: begin bcd3<=9;bcd2<=9;bcd1<=6;bcd0<=7; end
			9968: begin bcd3<=9;bcd2<=9;bcd1<=6;bcd0<=8; end
			9969: begin bcd3<=9;bcd2<=9;bcd1<=6;bcd0<=9; end
			9970: begin bcd3<=9;bcd2<=9;bcd1<=7;bcd0<=0; end
			9971: begin bcd3<=9;bcd2<=9;bcd1<=7;bcd0<=1; end
			9972: begin bcd3<=9;bcd2<=9;bcd1<=7;bcd0<=2; end
			9973: begin bcd3<=9;bcd2<=9;bcd1<=7;bcd0<=3; end
			9974: begin bcd3<=9;bcd2<=9;bcd1<=7;bcd0<=4; end
			9975: begin bcd3<=9;bcd2<=9;bcd1<=7;bcd0<=5; end
			9976: begin bcd3<=9;bcd2<=9;bcd1<=7;bcd0<=6; end
			9977: begin bcd3<=9;bcd2<=9;bcd1<=7;bcd0<=7; end
			9978: begin bcd3<=9;bcd2<=9;bcd1<=7;bcd0<=8; end
			9979: begin bcd3<=9;bcd2<=9;bcd1<=7;bcd0<=9; end
			9980: begin bcd3<=9;bcd2<=9;bcd1<=8;bcd0<=0; end
			9981: begin bcd3<=9;bcd2<=9;bcd1<=8;bcd0<=1; end
			9982: begin bcd3<=9;bcd2<=9;bcd1<=8;bcd0<=2; end
			9983: begin bcd3<=9;bcd2<=9;bcd1<=8;bcd0<=3; end
			9984: begin bcd3<=9;bcd2<=9;bcd1<=8;bcd0<=4; end
			9985: begin bcd3<=9;bcd2<=9;bcd1<=8;bcd0<=5; end
			9986: begin bcd3<=9;bcd2<=9;bcd1<=8;bcd0<=6; end
			9987: begin bcd3<=9;bcd2<=9;bcd1<=8;bcd0<=7; end
			9988: begin bcd3<=9;bcd2<=9;bcd1<=8;bcd0<=8; end
			9989: begin bcd3<=9;bcd2<=9;bcd1<=8;bcd0<=9; end
			9990: begin bcd3<=9;bcd2<=9;bcd1<=9;bcd0<=0; end
			9991: begin bcd3<=9;bcd2<=9;bcd1<=9;bcd0<=1; end
			9992: begin bcd3<=9;bcd2<=9;bcd1<=9;bcd0<=2; end
			9993: begin bcd3<=9;bcd2<=9;bcd1<=9;bcd0<=3; end
			9994: begin bcd3<=9;bcd2<=9;bcd1<=9;bcd0<=4; end
			9995: begin bcd3<=9;bcd2<=9;bcd1<=9;bcd0<=5; end
			9996: begin bcd3<=9;bcd2<=9;bcd1<=9;bcd0<=6; end
			9997: begin bcd3<=9;bcd2<=9;bcd1<=9;bcd0<=7; end
			9998: begin bcd3<=9;bcd2<=9;bcd1<=9;bcd0<=8; end
			9999: begin bcd3<=9;bcd2<=9;bcd1<=9;bcd0<=9; end

    endcase
    end
 
endmodule
